
module boothmul_Nbit16_DW01_inc_5 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] ;
  assign \carry[11]  = A[10];

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(\carry[11] ), .CO(\carry[12] ), .S(SUM[11]) );
  INV_X1 U1 ( .A(\carry[11] ), .ZN(SUM[10]) );
  XOR2_X1 U2 ( .A(\carry[31] ), .B(A[31]), .Z(SUM[31]) );
endmodule


module boothmul_Nbit16_DW01_inc_4 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ;
  assign \carry[12]  = A[11];

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  INV_X1 U1 ( .A(\carry[12] ), .ZN(SUM[11]) );
  XOR2_X1 U2 ( .A(\carry[31] ), .B(A[31]), .Z(SUM[31]) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n1) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U4 ( .A(n4), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n6), .A2(Ci), .ZN(n4) );
  XOR2_X1 U5 ( .A(A), .B(B), .Z(n6) );
  XOR2_X1 U6 ( .A(A), .B(B), .Z(n5) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n8), .Z(S) );
  NAND2_X1 U1 ( .A1(n5), .A2(n6), .ZN(n8) );
  NAND2_X1 U2 ( .A1(A), .A2(n4), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n1), .A2(B), .ZN(n6) );
  INV_X1 U5 ( .A(A), .ZN(n1) );
  INV_X1 U6 ( .A(B), .ZN(n4) );
  INV_X1 U7 ( .A(n7), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  NAND2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n1) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(n7), .ZN(Co) );
  XOR2_X1 U7 ( .A(A), .B(B), .Z(n8) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(n5), .A2(Ci), .ZN(n4) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  INV_X1 U1 ( .A(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n1), .A2(n8), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U7 ( .A(n8), .ZN(n4) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  INV_X2 U1 ( .A(n4), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  XOR2_X2 U4 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U5 ( .A(A), .B(B), .Z(n1) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  XOR2_X2 U1 ( .A(A), .B(B), .Z(n5) );
  INV_X2 U2 ( .A(n4), .ZN(Co) );
  AOI22_X2 U4 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(n5), .Z(n1) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X2 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X2 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n5), .A2(Ci), .ZN(n4) );
  XOR2_X1 U5 ( .A(A), .B(B), .Z(n5) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n5), .A2(Ci), .ZN(n4) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  XNOR2_X1 U1 ( .A(n4), .B(B), .ZN(n6) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n1) );
  INV_X1 U4 ( .A(A), .ZN(n4) );
  INV_X1 U5 ( .A(n5), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  XNOR2_X2 U2 ( .A(n1), .B(B), .ZN(n5) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(Co) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(B), .ZN(n5) );
  INV_X1 U4 ( .A(n4), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(n6), .A2(n7), .ZN(S) );
  NAND2_X1 U2 ( .A1(n4), .A2(n9), .ZN(n7) );
  INV_X1 U3 ( .A(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n5), .ZN(n6) );
  INV_X1 U6 ( .A(n8), .ZN(Co) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n1) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n9), .B2(n1), .ZN(n8) );
  INV_X1 U9 ( .A(n9), .ZN(n5) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  INV_X2 U1 ( .A(n5), .ZN(Co) );
  AOI22_X4 U2 ( .A1(n4), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
  XOR2_X2 U4 ( .A(B), .B(A), .Z(n6) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n1) );
  CLKBUF_X1 U6 ( .A(B), .Z(n4) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
  XOR2_X1 U2 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U3 ( .A(n1), .ZN(Co) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U1 ( .A(Ci), .B(n5), .Z(S) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n1) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(n1), .ZN(n4) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n1) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U4 ( .A(n4), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(n3), .B(Ci), .Z(S) );
  XOR2_X2 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(n5), .A2(Ci), .ZN(n4) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  INV_X2 U1 ( .A(n4), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  XNOR2_X2 U4 ( .A(n1), .B(B), .ZN(n5) );
  INV_X1 U5 ( .A(A), .ZN(n1) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Co) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(Ci), .B(n3), .Z(S) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  XNOR2_X1 U1 ( .A(n4), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(A), .ZN(n4) );
  INV_X1 U5 ( .A(n5), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  NAND2_X2 U1 ( .A1(n4), .A2(n3), .ZN(Co) );
  XNOR2_X2 U2 ( .A(n5), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(A), .ZN(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U6 ( .A1(n6), .A2(Ci), .ZN(n4) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n8), .Z(S) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
  NAND2_X1 U2 ( .A1(A), .A2(n4), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n1), .A2(B), .ZN(n6) );
  NAND2_X2 U5 ( .A1(n5), .A2(n6), .ZN(n8) );
  INV_X1 U6 ( .A(A), .ZN(n1) );
  INV_X1 U7 ( .A(B), .ZN(n4) );
  INV_X1 U8 ( .A(n7), .ZN(Co) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  INV_X1 U1 ( .A(n8), .ZN(n4) );
  INV_X1 U2 ( .A(n7), .ZN(Co) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n1), .A2(n8), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(S) );
  INV_X1 U7 ( .A(Ci), .ZN(n1) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U3 ( .A(n6), .B(Ci), .Z(S) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U4 ( .A1(n6), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
  INV_X1 U6 ( .A(A), .ZN(n5) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U1 ( .A1(n5), .A2(Ci), .ZN(n4) );
  NAND2_X1 U2 ( .A1(n4), .A2(n3), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n1) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n6) );
  INV_X1 U4 ( .A(n5), .ZN(Co) );
  AOI22_X1 U5 ( .A1(n4), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(B), .Z(n4) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8, n9;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U1 ( .A1(n6), .A2(n7), .ZN(S) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n5), .ZN(n6) );
  INV_X1 U3 ( .A(n8), .ZN(Co) );
  CLKBUF_X1 U5 ( .A(Ci), .Z(n1) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n9), .B2(n1), .ZN(n8) );
  NAND2_X1 U7 ( .A1(n4), .A2(n9), .ZN(n7) );
  INV_X1 U8 ( .A(Ci), .ZN(n4) );
  INV_X1 U9 ( .A(n9), .ZN(n5) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7;

  NAND2_X2 U1 ( .A1(n7), .A2(Ci), .ZN(n5) );
  NAND2_X2 U2 ( .A1(n4), .A2(n5), .ZN(Co) );
  XOR2_X2 U3 ( .A(Ci), .B(n1), .Z(S) );
  CLKBUF_X1 U4 ( .A(n7), .Z(n1) );
  XOR2_X1 U5 ( .A(A), .B(B), .Z(n7) );
  NAND2_X1 U6 ( .A1(n6), .A2(A), .ZN(n4) );
  CLKBUF_X1 U7 ( .A(B), .Z(n6) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U1 ( .A(Ci), .B(n5), .Z(S) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n1) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(n1), .ZN(n4) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n1) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U4 ( .A(n4), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X2 U1 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(Co) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(n5), .A2(Ci), .ZN(n4) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  INV_X1 U1 ( .A(n7), .ZN(Co) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n1), .A2(n8), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U6 ( .A(Ci), .ZN(n1) );
  INV_X1 U7 ( .A(n8), .ZN(n4) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  AOI22_X4 U1 ( .A1(n1), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  INV_X2 U2 ( .A(n4), .ZN(Co) );
  XOR2_X2 U4 ( .A(B), .B(A), .Z(n5) );
  CLKBUF_X1 U5 ( .A(B), .Z(n1) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X2 U1 ( .A(n1), .ZN(Co) );
  AOI22_X4 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  NAND2_X2 U1 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n6), .ZN(S) );
  INV_X1 U3 ( .A(n7), .ZN(Co) );
  INV_X1 U5 ( .A(Ci), .ZN(n1) );
  NAND2_X1 U6 ( .A1(n1), .A2(n8), .ZN(n6) );
  INV_X1 U7 ( .A(n8), .ZN(n4) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  INV_X2 U1 ( .A(n5), .ZN(Co) );
  NOR2_X4 U2 ( .A1(n1), .A2(n4), .ZN(n5) );
  AND2_X4 U4 ( .A1(n6), .A2(Ci), .ZN(n4) );
  AND2_X1 U5 ( .A1(B), .A2(A), .ZN(n1) );
  XOR2_X2 U6 ( .A(A), .B(B), .Z(n6) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n5), .B(Ci), .Z(S) );
  INV_X1 U1 ( .A(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(B), .ZN(n5) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(Co) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XNOR2_X1 U1 ( .A(n1), .B(B), .ZN(n5) );
  INV_X1 U2 ( .A(A), .ZN(n1) );
  INV_X1 U4 ( .A(n4), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X1 U1 ( .A1(n5), .A2(Ci), .ZN(n4) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XNOR2_X1 U1 ( .A(B), .B(n5), .ZN(n6) );
  AND2_X1 U2 ( .A1(n6), .A2(Ci), .ZN(n4) );
  OR2_X1 U4 ( .A1(n3), .A2(n4), .ZN(Co) );
  AND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
  INV_X1 U6 ( .A(A), .ZN(n5) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  NAND2_X1 U1 ( .A1(n5), .A2(n6), .ZN(S) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n8) );
  INV_X1 U4 ( .A(n8), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n1), .A2(n8), .ZN(n6) );
  INV_X1 U6 ( .A(Ci), .ZN(n1) );
  INV_X1 U7 ( .A(n7), .ZN(Co) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U1 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U1 ( .A1(n5), .A2(Ci), .ZN(n4) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U1 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
  AOI22_X1 U3 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n1), .Z(S) );
  XNOR2_X1 U1 ( .A(n4), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n4), .B(B), .ZN(n6) );
  INV_X1 U4 ( .A(A), .ZN(n4) );
  INV_X1 U5 ( .A(n5), .ZN(Co) );
  AOI22_X1 U6 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U1 ( .A1(n5), .A2(n6), .ZN(S) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(n5) );
  INV_X1 U3 ( .A(n8), .ZN(n4) );
  INV_X1 U5 ( .A(n7), .ZN(Co) );
  NAND2_X1 U6 ( .A1(n1), .A2(n8), .ZN(n6) );
  INV_X1 U7 ( .A(Ci), .ZN(n1) );
  AOI22_X1 U8 ( .A1(B), .A2(A), .B1(n8), .B2(Ci), .ZN(n7) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  INV_X1 U1 ( .A(n6), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n4) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
  INV_X1 U6 ( .A(n5), .ZN(Co) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U4 ( .A(n1), .ZN(Co) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n1) );
  INV_X1 U2 ( .A(n5), .ZN(Co) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n1), .B2(n4), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n4) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  INV_X2 U1 ( .A(n4), .ZN(Co) );
  AOI22_X2 U2 ( .A1(n1), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n5) );
  XOR2_X1 U4 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U5 ( .A(B), .Z(n1) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6, n7, n8;

  XOR2_X1 U3 ( .A(Ci), .B(n8), .Z(S) );
  NAND2_X1 U1 ( .A1(A), .A2(n4), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n1), .A2(B), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(n8) );
  INV_X1 U5 ( .A(A), .ZN(n1) );
  INV_X1 U6 ( .A(B), .ZN(n4) );
  AOI22_X2 U7 ( .A1(B), .A2(A), .B1(Ci), .B2(n8), .ZN(n7) );
  INV_X1 U8 ( .A(n7), .ZN(Co) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n1), .B2(Ci), .ZN(n4) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U5 ( .A1(n5), .A2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X2 U1 ( .A(A), .B(B), .Z(n3) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U4 ( .A(n1), .ZN(Co) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Co) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n6), .Z(S) );
  NAND2_X2 U1 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(n6), .A2(Ci), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n5), .A2(A), .ZN(n4) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n6) );
  CLKBUF_X1 U6 ( .A(B), .Z(n5) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(Ci), .B2(n3), .ZN(n1) );
  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(Co) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(n4) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  INV_X1 U1 ( .A(n1), .ZN(Co) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n3) );
  XOR2_X1 U3 ( .A(n3), .B(Ci), .Z(S) );
  AOI22_X1 U4 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  INV_X2 U1 ( .A(n5), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n6), .B2(Ci), .ZN(n5) );
  XOR2_X2 U4 ( .A(A), .B(B), .Z(n6) );
  INV_X1 U5 ( .A(n6), .ZN(n1) );
  INV_X1 U6 ( .A(n1), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  NAND2_X2 U1 ( .A1(n5), .A2(Ci), .ZN(n4) );
  NAND2_X2 U2 ( .A1(n4), .A2(n3), .ZN(Co) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n3) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI22_X2 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n1) );
  XOR2_X2 U4 ( .A(A), .B(B), .Z(n3) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n1), .B2(Ci), .ZN(n4) );
endmodule


module MUX21_GENERIC_N4_55 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_55 UIV ( .A(SEL), .Y(SB) );
  ND2_660 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_659 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_658 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_657 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_656 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_655 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_654 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_653 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_652 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_651 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_650 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_649 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_54 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_54 UIV ( .A(SEL), .Y(SB) );
  ND2_648 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_647 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_646 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_645 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_644 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_643 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_642 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_641 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_640 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_639 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_638 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_637 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_53 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_53 UIV ( .A(SEL), .Y(SB) );
  ND2_636 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_635 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_634 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_633 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_632 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_631 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_630 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_629 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_628 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_627 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_626 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_625 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_52 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_52 UIV ( .A(SEL), .Y(SB) );
  ND2_624 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_623 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_622 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_621 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_620 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_619 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_618 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_617 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_616 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_615 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_614 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_613 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_51 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_51 UIV ( .A(SEL), .Y(SB) );
  ND2_612 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_611 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_610 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_609 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_608 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_607 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_606 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_605 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_604 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_603 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_602 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_601 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_50 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_50 UIV ( .A(SEL), .Y(SB) );
  ND2_600 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_599 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_598 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_597 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_596 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_595 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_594 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_593 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_592 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_591 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_590 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_589 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_49 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_49 UIV ( .A(SEL), .Y(SB) );
  ND2_588 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_587 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_586 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_585 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_584 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_583 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_582 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_581 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_580 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_579 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_578 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_577 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_48 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_48 UIV ( .A(SEL), .Y(SB) );
  ND2_576 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_575 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_574 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_573 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_572 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_571 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_570 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_569 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_568 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_567 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_566 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_565 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_47 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_47 UIV ( .A(SEL), .Y(SB) );
  ND2_564 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_563 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_562 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_561 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_560 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_559 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_558 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_557 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_556 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_555 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_554 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_553 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_46 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_46 UIV ( .A(SEL), .Y(SB) );
  ND2_552 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_551 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_550 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_549 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_548 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_547 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_546 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_545 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_544 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_543 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_542 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_541 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_45 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_45 UIV ( .A(SEL), .Y(SB) );
  ND2_540 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_539 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_538 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_537 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_536 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_535 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_534 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_533 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_532 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_531 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_530 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_529 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_44 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB, n1;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_44 UIV ( .A(SEL), .Y(SB) );
  ND2_528 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_527 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_526 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_525 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_524 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_523 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_522 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_521 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_520 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_519 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_518 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_517 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  CLKBUF_X1 U1 ( .A(SEL), .Z(n1) );
endmodule


module MUX21_GENERIC_N4_43 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_43 UIV ( .A(SEL), .Y(SB) );
  ND2_516 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_515 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_514 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_513 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_512 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_511 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_510 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_509 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_508 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_507 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_506 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_505 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_42 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_42 UIV ( .A(SEL), .Y(SB) );
  ND2_504 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_503 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_502 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_501 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_500 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_499 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_498 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_497 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_496 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_495 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_494 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_493 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_41 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_41 UIV ( .A(SEL), .Y(SB) );
  ND2_492 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_491 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_490 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_489 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_488 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_487 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_486 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_485 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_484 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_483 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_482 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_481 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_40 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_40 UIV ( .A(SEL), .Y(SB) );
  ND2_480 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_479 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_478 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_477 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_476 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_475 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_474 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_473 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_472 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_471 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_470 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_469 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_39 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_39 UIV ( .A(SEL), .Y(SB) );
  ND2_468 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_467 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_466 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_465 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_464 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_463 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_462 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_461 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_460 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_459 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_458 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_457 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_38 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_38 UIV ( .A(SEL), .Y(SB) );
  ND2_456 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_455 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_454 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_453 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_452 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_451 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_450 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_449 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_448 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_447 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_446 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_445 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_37 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_37 UIV ( .A(SEL), .Y(SB) );
  ND2_444 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_443 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_442 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_441 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_440 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_439 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_438 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_437 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_436 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_435 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_434 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_433 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_36 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_36 UIV ( .A(SEL), .Y(SB) );
  ND2_432 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_431 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_430 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_429 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_428 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_427 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_426 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_425 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_424 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_423 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_422 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_421 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_35 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_35 UIV ( .A(SEL), .Y(SB) );
  ND2_420 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_419 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_418 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_417 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_416 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_415 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_414 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_413 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_412 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_411 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_410 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_409 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_34 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_34 UIV ( .A(SEL), .Y(SB) );
  ND2_408 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_407 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_406 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_405 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_404 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_403 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_402 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_401 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_400 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_399 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_398 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_397 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_33 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_33 UIV ( .A(SEL), .Y(SB) );
  ND2_396 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_395 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_394 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_393 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_392 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_391 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_390 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_389 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_388 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_387 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_386 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_385 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_32 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_32 UIV ( .A(SEL), .Y(SB) );
  ND2_384 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_383 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_382 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_381 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_380 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_379 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_378 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_377 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_376 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_375 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_374 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_373 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_31 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_31 UIV ( .A(SEL), .Y(SB) );
  ND2_372 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_371 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_370 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_369 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_368 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_367 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_366 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_365 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_364 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_363 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_362 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_361 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_30 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_30 UIV ( .A(SEL), .Y(SB) );
  ND2_360 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_359 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_358 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_357 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_356 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_355 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_354 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_353 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_352 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_351 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_350 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_349 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_29 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_29 UIV ( .A(SEL), .Y(SB) );
  ND2_348 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_347 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_346 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_345 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_344 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_343 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_342 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_341 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_340 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_339 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_338 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_337 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_28 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_28 UIV ( .A(SEL), .Y(SB) );
  ND2_336 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_335 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_334 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_333 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_332 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_331 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_330 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_329 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_328 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_327 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_326 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_325 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_27 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_27 UIV ( .A(SEL), .Y(SB) );
  ND2_324 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_323 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_322 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_321 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_320 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_319 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_318 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_317 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_316 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_315 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_314 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_313 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_26 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_26 UIV ( .A(SEL), .Y(SB) );
  ND2_312 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_311 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_310 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_309 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_308 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_307 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_306 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_305 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_304 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_303 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_302 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_301 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_25 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_25 UIV ( .A(SEL), .Y(SB) );
  ND2_300 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_299 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_298 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_297 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_296 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_295 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_294 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_293 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_292 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_291 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_290 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_289 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_24 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_24 UIV ( .A(SEL), .Y(SB) );
  ND2_288 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_287 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_286 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_285 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_284 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_283 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_282 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_281 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_280 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_279 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_278 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_277 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_23 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_23 UIV ( .A(SEL), .Y(SB) );
  ND2_276 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_275 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_274 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_273 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_272 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_271 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_270 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_269 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_268 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_267 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_266 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_265 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_22 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_22 UIV ( .A(SEL), .Y(SB) );
  ND2_264 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_263 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_262 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_261 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_260 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_259 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_258 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_257 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_256 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_255 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_254 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_253 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_21 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_21 UIV ( .A(SEL), .Y(SB) );
  ND2_252 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_251 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_250 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_249 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_248 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_247 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_246 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_245 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_244 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_243 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_242 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_241 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_20 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_20 UIV ( .A(SEL), .Y(SB) );
  ND2_240 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_239 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_238 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_237 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_236 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_235 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_234 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_233 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_232 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_231 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_230 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_229 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_19 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_19 UIV ( .A(SEL), .Y(SB) );
  ND2_228 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_227 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_226 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_225 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_224 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_223 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_222 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_221 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_220 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_219 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_218 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_217 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_18 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_18 UIV ( .A(SEL), .Y(SB) );
  ND2_216 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_215 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_214 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_213 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_212 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_211 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_210 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_209 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_208 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_207 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_206 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_205 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_17 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_17 UIV ( .A(SEL), .Y(SB) );
  ND2_204 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_203 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_202 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_201 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_200 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_199 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_198 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_197 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_196 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_195 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_194 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_193 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_16 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_16 UIV ( .A(SEL), .Y(SB) );
  ND2_192 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_191 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_190 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_189 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_188 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_187 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_186 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_185 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_184 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_183 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_182 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_181 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_15 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_15 UIV ( .A(SEL), .Y(SB) );
  ND2_180 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_179 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_178 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_177 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_176 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_175 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_174 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_173 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_172 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_171 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_170 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_169 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_14 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_14 UIV ( .A(SEL), .Y(SB) );
  ND2_168 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_167 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_166 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_165 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_164 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_163 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_162 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_161 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_160 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_159 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_158 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_157 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_13 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_13 UIV ( .A(SEL), .Y(SB) );
  ND2_156 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_155 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_154 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_153 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_152 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_151 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_150 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_149 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_148 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_147 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_146 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_145 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_12 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_12 UIV ( .A(SEL), .Y(SB) );
  ND2_144 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_143 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_142 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_141 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_140 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_139 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_138 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_137 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_136 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_135 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_134 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_133 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_11 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_11 UIV ( .A(SEL), .Y(SB) );
  ND2_132 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_131 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_130 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_129 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_128 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_127 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_126 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_125 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_124 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_123 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_122 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_121 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_10 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_10 UIV ( .A(SEL), .Y(SB) );
  ND2_120 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_119 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_118 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_117 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_116 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_115 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_114 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_113 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_112 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_111 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_110 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_109 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_9 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_9 UIV ( .A(SEL), .Y(SB) );
  ND2_108 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_107 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_106 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_105 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_104 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_103 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_102 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_101 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_100 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_99 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_98 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_97 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_8 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_8 UIV ( .A(SEL), .Y(SB) );
  ND2_96 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_95 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_94 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_93 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_92 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_91 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_90 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_89 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_88 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_87 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_86 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_85 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_7 UIV ( .A(SEL), .Y(SB) );
  ND2_84 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_83 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_82 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_81 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_80 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_79 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_78 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_77 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_76 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_75 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_74 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_73 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_6 UIV ( .A(SEL), .Y(SB) );
  ND2_72 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_71 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_70 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_69 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_68 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_67 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_66 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_65 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_64 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_63 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_62 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_61 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_5 UIV ( .A(SEL), .Y(SB) );
  ND2_60 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_59 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_58 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_57 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_56 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_55 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_54 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_53 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_52 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_51 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_50 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_49 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_4 UIV ( .A(SEL), .Y(SB) );
  ND2_48 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_47 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_46 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_45 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_44 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_43 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_42 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_41 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_40 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_39 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_38 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_37 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_3 UIV ( .A(SEL), .Y(SB) );
  ND2_36 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_35 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_34 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_33 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_32 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_31 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_30 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_29 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_28 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_27 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_26 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_25 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_2 UIV ( .A(SEL), .Y(SB) );
  ND2_24 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_23 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_22 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_21 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_20 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_19 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_18 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_17 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_16 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_15 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_14 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_13 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_1 UIV ( .A(SEL), .Y(SB) );
  ND2_12 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_11 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_10 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_9 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_8 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_7 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_6 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_5 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_4 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_2 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_1 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module RCA_generic_N4_111 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_444 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_443 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_442 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_441 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_110 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_440 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_439 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_438 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_437 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_109 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_436 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_435 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_434 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_433 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_108 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_432 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_431 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_430 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_429 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_107 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_428 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_427 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_426 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_425 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_106 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_424 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_423 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_422 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_421 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_105 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_420 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_419 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_418 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_417 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_104 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_416 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_415 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_414 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_413 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_103 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_412 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_411 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_410 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_409 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_102 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_408 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_407 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_406 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_405 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_101 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_404 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_403 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_402 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_401 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_100 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_400 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_399 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_398 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_397 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_99 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_396 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_395 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_394 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_393 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_98 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_392 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_391 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_390 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_389 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_97 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_388 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_387 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_386 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_385 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_96 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_384 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_383 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_382 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_381 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_95 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_380 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_379 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_378 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_377 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_94 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_376 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_375 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_374 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_373 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_93 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_372 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_371 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_370 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_369 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_92 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_368 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_367 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_366 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_365 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_91 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_364 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_363 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_362 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_361 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_90 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_360 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_359 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_358 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_357 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_89 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_356 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_355 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_354 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_353 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_88 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_352 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_351 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_350 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_349 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_87 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_348 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_347 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_346 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_345 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_86 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_344 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_343 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_342 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_341 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_85 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_340 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_339 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_338 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_337 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_84 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_336 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_335 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_334 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_333 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_83 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_332 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_331 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_330 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_329 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_82 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_328 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_327 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_326 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_325 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_81 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_324 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_323 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_322 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_321 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_80 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_320 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_319 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_318 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_317 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_79 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_316 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_315 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_314 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_313 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_78 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_312 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_311 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_310 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_309 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_77 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_308 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_307 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_306 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_305 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_76 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_304 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_303 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_302 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_301 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_75 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_300 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_299 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_298 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_297 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_74 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_296 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_295 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_294 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_293 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_73 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_292 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_291 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_290 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_289 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_72 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_288 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_287 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_286 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_285 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_71 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_284 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_283 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_282 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_281 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_70 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_280 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_279 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_278 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_277 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_69 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_276 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_275 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_274 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_273 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_68 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_272 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_271 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_270 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_269 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_67 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_268 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_267 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_266 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_265 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_66 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_264 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_263 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_262 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_261 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_65 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_260 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_259 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_258 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_257 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_64 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_256 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_255 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_254 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_253 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_63 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_252 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_251 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_250 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_249 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_248 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_247 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_246 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_245 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_61 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_244 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_243 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_242 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_241 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_240 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_239 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_238 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_237 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_59 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_236 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_235 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_234 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_233 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_232 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_231 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_230 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_229 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_57 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_228 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_227 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_226 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_225 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_224 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_223 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_222 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_221 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_55 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_220 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_219 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_218 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_217 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_216 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_215 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_214 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_213 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_53 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_212 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_211 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_210 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_209 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_208 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_207 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_206 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_205 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_51 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_204 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_203 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_202 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_201 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_200 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_199 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_198 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_197 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_49 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_196 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_195 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_194 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_193 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_48 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_192 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_191 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_190 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_189 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_47 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_188 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_187 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_186 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_185 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_46 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_184 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_183 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_182 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_181 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_45 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_180 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_179 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_178 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_177 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_44 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_176 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_175 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_174 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_173 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_43 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_172 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_171 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_170 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_169 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_42 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_168 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_167 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_166 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_165 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_41 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_164 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_163 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_162 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_161 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_40 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_160 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_159 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_158 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_157 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_39 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_156 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_155 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_154 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_153 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_38 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_152 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_151 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_150 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_149 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_37 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_148 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_147 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_146 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_145 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_36 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_144 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_143 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_142 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_141 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_35 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_140 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_139 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_138 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_137 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_34 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_136 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_135 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_134 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_133 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_33 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_132 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_131 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_130 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_129 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_128 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_124 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_123 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_122 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_121 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_120 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_119 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_118 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_117 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_116 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_115 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_114 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_113 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_108 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_107 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_106 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_105 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_104 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_103 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_102 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_101 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_100 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_99 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_98 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_97 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_96 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_95 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_92 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_91 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_90 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_89 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_88 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_87 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_86 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_85 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_84 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_83 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_82 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_81 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_80 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_79 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_78 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_77 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_76 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_75 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_74 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_73 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_72 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_71 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_70 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_69 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_68 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_67 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_66 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_65 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module cs_generic_N4_55 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_110 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_109 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_55 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_54 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_108 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_107 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_54 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_53 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_106 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_105 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_53 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_52 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_104 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_103 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_52 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_51 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_102 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_101 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_51 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_50 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_100 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_99 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_50 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_49 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_98 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_97 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_49 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_48 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_96 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_95 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_48 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_47 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_94 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_93 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_47 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_46 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_92 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_91 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_46 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_45 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_90 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_89 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_45 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_44 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_88 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_87 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_44 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_43 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_86 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_85 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_43 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_42 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_84 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_83 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_42 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_41 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_82 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_81 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_41 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_40 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_80 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_79 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_40 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_39 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_78 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_77 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_39 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_38 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_76 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_75 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_38 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_37 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_74 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_73 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_37 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_36 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_72 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_71 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_36 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_35 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_70 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_69 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_35 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_34 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_68 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_67 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_34 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_33 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_66 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_65 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_33 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_32 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_64 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_63 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_32 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_31 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_62 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_61 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_31 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_30 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_60 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_59 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_30 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_29 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_58 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_57 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_29 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_28 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_56 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_55 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_28 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_27 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_54 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_53 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_27 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_26 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_52 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_51 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_26 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_25 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_50 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_49 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_25 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_24 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_48 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_47 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_24 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_23 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_46 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_45 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_23 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_22 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_44 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_43 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_22 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_21 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_42 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_41 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_21 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_20 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_40 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_39 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_20 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_19 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_38 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_37 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_19 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_18 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_36 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_35 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_18 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_17 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_34 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_33 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_17 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_16 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_32 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_31 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_16 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_30 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_29 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_15 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_28 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_27 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_14 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_26 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_25 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_13 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_24 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_23 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_12 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_22 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_21 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_11 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_20 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_19 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_10 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_18 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_17 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_9 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_16 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_15 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_8 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_14 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_13 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_7 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_12 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_11 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_6 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_10 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_9 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_5 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_8 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_7 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_4 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_6 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_5 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_3 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_4 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_3 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_2 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_2 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_1 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_1 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module block_pg_188 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_187 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_186 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_185 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_184 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_183 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_182 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_181 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X2 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_pg_180 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_179 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_178 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_177 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_176 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_175 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_174 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_173 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_172 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X2 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_171 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X2 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_170 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_169 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_168 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_167 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_166 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_165 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_164 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_163 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_162 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_161 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_160 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_159 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_158 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_157 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_156 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_155 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_154 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_153 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_152 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_151 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_150 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_149 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_148 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_147 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_146 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_145 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_144 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X2 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_143 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_142 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_141 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_140 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_139 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_138 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_137 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_136 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_135 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_134 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_133 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_132 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_131 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_130 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_129 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_128 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_127 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X2 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X2 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_126 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_125 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pik), .A2(Pk1j), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_124 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_123 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_122 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_121 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_120 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_119 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_118 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_117 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_116 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X2 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_115 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_114 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_113 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_112 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X2 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_111 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_110 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_109 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_108 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_107 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_106 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_105 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_104 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_103 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_102 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_101 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_100 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_99 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_98 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X2 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_97 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_96 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_95 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_94 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_93 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_92 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_91 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_90 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_89 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_88 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AND2_X2 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X2 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_87 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_86 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_85 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_84 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_83 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_82 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_81 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_80 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_79 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_78 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_77 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_76 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_75 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_74 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_73 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pik), .A2(Pk1j), .ZN(Pij) );
endmodule


module block_pg_72 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_71 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_70 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_69 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_68 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_67 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_66 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_65 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_64 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_63 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n2, n3, n4;

  OR2_X1 U1 ( .A1(n4), .A2(Gik), .ZN(Gij) );
  INV_X1 U2 ( .A(Pik), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n2), .A2(n3), .ZN(n4) );
  INV_X1 U4 ( .A(Gk1j), .ZN(n2) );
  AND2_X1 U5 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_62 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_61 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AND2_X2 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X2 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_60 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_59 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_58 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_57 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_56 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_55 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X2 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X2 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_54 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_53 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_52 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_51 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_50 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_49 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_48 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_47 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_46 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_45 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_44 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_43 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_42 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  AND2_X2 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_41 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_40 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_39 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_38 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_37 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_36 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_35 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(n2), .A2(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U3 ( .A1(Gk1j), .A2(Pik), .ZN(n2) );
  INV_X1 U4 ( .A(Gik), .ZN(n3) );
endmodule


module block_pg_34 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AND2_X2 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X2 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_33 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_32 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_31 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_30 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_29 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_28 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_27 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_26 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_25 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_24 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_23 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_22 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_21 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_20 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_19 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_18 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_17 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Gij) );
endmodule


module block_pg_16 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_15 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_14 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_13 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_12 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_11 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_10 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_9 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_8 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(n2), .A2(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  NAND2_X1 U3 ( .A1(Gk1j), .A2(Pik), .ZN(n2) );
  INV_X1 U4 ( .A(Gik), .ZN(n3) );
endmodule


module block_pg_7 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_6 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_5 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_4 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_3 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_2 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
endmodule


module block_pg_1 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_g_69 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_68 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_67 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_66 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_65 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_64 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_63 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_62 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_61 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X4 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X4 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_60 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_59 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_58 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_57 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_56 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X4 U2 ( .A(n1), .ZN(Gij) );
endmodule


module block_g_55 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_54 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_53 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_52 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X4 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X4 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_51 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_50 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_49 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_48 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_47 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_46 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_45 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_44 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_43 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_42 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X4 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X4 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_41 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_40 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_39 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_38 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_37 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_36 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X2 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_35 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_34 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_33 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Gij) );
endmodule


module block_g_32 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Gij) );
endmodule


module block_g_31 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_30 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_29 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_28 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_27 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_26 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_25 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_24 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_23 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Gij) );
endmodule


module block_g_22 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_21 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Gij) );
endmodule


module block_g_20 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_19 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_18 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_17 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_16 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X2 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_15 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_14 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_13 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  AOI21_X2 U1 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Gij) );
endmodule


module block_g_12 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2, n3, n4;

  OR2_X4 U1 ( .A1(n4), .A2(Gik), .ZN(Gij) );
  NOR2_X2 U2 ( .A1(n2), .A2(n3), .ZN(n4) );
  INV_X1 U3 ( .A(Pik), .ZN(n2) );
  INV_X1 U4 ( .A(Gk1j), .ZN(n3) );
endmodule


module block_g_11 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_10 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_9 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_8 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_7 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_6 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_5 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_4 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_3 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_2 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module block_g_1 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n1) );
endmodule


module ND2_3743 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3742 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3741 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3740 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3739 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3738 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3737 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3736 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3735 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3734 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3733 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3732 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3731 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3730 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3729 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3728 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3727 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3726 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3725 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3724 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3723 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3722 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3721 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3720 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3719 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3718 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3717 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3716 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3715 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3714 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3713 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3712 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3711 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3710 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3709 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3708 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3707 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3706 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3705 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3704 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3703 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3702 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3701 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3700 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3699 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3698 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3697 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_3696 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3695 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3694 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_3693 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3692 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3691 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3690 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3689 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3688 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3687 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3686 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3685 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3684 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_3683 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3682 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_3681 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3680 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3679 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3678 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3677 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3676 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3675 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3674 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3673 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3672 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3671 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3670 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3669 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3668 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3667 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3666 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3665 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3664 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3663 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3662 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3661 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3660 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3659 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3658 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3657 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3656 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3655 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3654 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3653 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3652 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3651 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3650 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3649 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3648 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3647 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3646 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3645 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3644 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3643 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3642 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3641 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3640 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3639 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3638 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3637 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3636 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3635 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3634 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3633 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3632 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3631 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3630 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3629 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3628 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3627 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3626 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3625 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3624 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3623 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3622 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3621 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3620 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3619 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3618 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3617 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3616 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3615 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3614 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3613 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3612 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3611 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3610 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3609 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3608 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3607 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3606 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3605 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3604 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3603 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3602 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3601 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3600 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3599 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3598 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3597 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3596 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3595 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3594 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3593 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3592 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3591 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3590 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3589 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3588 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3587 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3586 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3585 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3584 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3583 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3582 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3581 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3580 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3579 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3578 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3577 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3576 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3575 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3574 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3573 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3572 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3571 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3570 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3569 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3568 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3567 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3566 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3565 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3564 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3563 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3562 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3561 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3560 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3559 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3558 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3557 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3556 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3555 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3554 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3553 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3552 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3551 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3550 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3549 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3548 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3547 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3546 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3545 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3544 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3543 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3542 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3541 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3540 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3539 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3538 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3537 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3536 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3535 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3534 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3533 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3532 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3531 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3530 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3529 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3528 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3527 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3526 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3525 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3524 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3523 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3522 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3521 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3520 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3519 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3518 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3517 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3516 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3515 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3514 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3513 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3512 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3511 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3510 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3509 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3508 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3507 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3506 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3505 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3504 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3503 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3502 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3501 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3500 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3499 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3498 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3497 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3496 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3495 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3494 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3493 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3492 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3491 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3490 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3489 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3488 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3487 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3486 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3485 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3484 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3483 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3482 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3481 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3480 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3479 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3478 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3477 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3476 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3475 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3474 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3473 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3472 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3471 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3470 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3469 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3468 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3467 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3466 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3465 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3464 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3463 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3462 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3461 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3460 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3459 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3458 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3457 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3456 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3455 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3454 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3453 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3452 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3451 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3450 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3449 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3448 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3447 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3446 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3445 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3444 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3443 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3442 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3441 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3440 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3439 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3438 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3437 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3436 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3435 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3434 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3433 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3432 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3431 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3430 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3429 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3428 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3427 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3426 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3425 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3424 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3423 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3422 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3421 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3420 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3419 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3418 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3417 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3416 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3415 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3414 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3413 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3412 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3411 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3410 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3409 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3408 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3407 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3406 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3405 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3404 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3403 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3402 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3401 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3400 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3399 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3398 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3397 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3396 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3395 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3394 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_3393 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3392 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3391 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3390 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3389 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3388 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3387 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3386 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3385 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3384 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3383 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3382 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3381 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3380 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3379 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3378 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3377 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3376 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3375 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3374 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3373 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3372 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3371 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3370 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3369 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3368 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3367 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3366 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3365 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3364 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3363 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3362 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3361 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3360 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3359 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3358 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3357 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3356 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3355 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3354 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3353 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3352 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3351 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3350 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3349 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3348 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3347 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3346 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3345 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3344 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3343 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3342 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3341 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3340 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3339 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3338 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3337 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3336 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3335 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3334 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3333 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3332 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3331 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3330 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3329 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3328 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3327 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3326 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3325 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3324 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3323 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3322 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3321 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3320 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3319 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3318 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3317 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3316 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3315 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_3314 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3313 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3312 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3311 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3310 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3309 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3308 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3307 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3306 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3305 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3304 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3303 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3302 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3301 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3300 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3299 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3298 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3297 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3296 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3295 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3294 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3293 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3292 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3291 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3290 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3289 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3288 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3287 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3286 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3285 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3284 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3283 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3282 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3281 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3280 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3279 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3278 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3277 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3276 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3275 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3274 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3273 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3272 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3271 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3270 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3269 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3268 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3267 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3266 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3265 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3264 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3263 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3262 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3261 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3260 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3259 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3258 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3257 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3256 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3255 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3254 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3253 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3252 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3251 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3250 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3249 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3248 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3247 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3246 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3245 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3244 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3243 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3242 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3241 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3240 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3239 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3238 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3237 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3236 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3235 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3234 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3233 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3232 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3231 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3230 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3229 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3228 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3227 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3226 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3225 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3224 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3223 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3222 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3221 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3220 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3219 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3218 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3217 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3216 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3215 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3214 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3213 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3212 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3211 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3210 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3209 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3208 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3207 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3206 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3205 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3204 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3203 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3202 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3201 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3200 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3199 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3198 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3197 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3196 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3195 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3194 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3193 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3192 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3191 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3190 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3189 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3188 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3187 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3186 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3185 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3184 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3183 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3182 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3181 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3180 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3179 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3178 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3177 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3176 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3175 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3174 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3173 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3172 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3171 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3170 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3169 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3168 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3167 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3166 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3165 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3164 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3163 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3162 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3161 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3160 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3159 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3158 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3157 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3156 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3155 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3154 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3153 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3152 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3151 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3150 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3149 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3148 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3147 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3146 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3145 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3144 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3143 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3142 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3141 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3140 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3139 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3138 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3137 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3136 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3135 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3134 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3133 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3132 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3131 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3130 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3129 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3128 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3127 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3126 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3125 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3124 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3123 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3122 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3121 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3120 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3119 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3118 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3117 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3116 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3115 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3114 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3113 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3112 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3111 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3110 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3109 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3108 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3107 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3106 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3105 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3104 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3103 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3102 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3101 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3100 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3099 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3098 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3097 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3096 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3095 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3094 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3093 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3092 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3091 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3090 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3089 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3088 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3087 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3086 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3085 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3084 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3083 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3082 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3081 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3080 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3079 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3078 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3077 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3076 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3075 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3074 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3073 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3072 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3071 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3070 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3069 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3068 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3067 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3066 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3065 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3064 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3063 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3062 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3061 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3060 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3059 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3058 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3057 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3056 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3055 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3054 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3053 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3052 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3051 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3050 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3049 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3048 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3047 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3046 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3045 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3044 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3043 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3042 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3041 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3040 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3039 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3038 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3037 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3036 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3035 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3034 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3033 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3032 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3031 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3030 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3029 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3028 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3027 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3026 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3025 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3024 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3023 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3022 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3021 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3020 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3019 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3018 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3017 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3016 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3015 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3014 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3013 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3012 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3011 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3010 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3009 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3008 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3007 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3006 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3005 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3004 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3003 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3002 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3001 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3000 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2999 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2998 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2997 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2996 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2995 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2994 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2993 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2992 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2991 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2990 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2989 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2988 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2987 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2986 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2985 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2984 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2983 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2982 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2981 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2980 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2979 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2978 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2977 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2976 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2975 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2974 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2973 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2972 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2971 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2970 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2969 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2968 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2967 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2966 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2965 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2964 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2963 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2962 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2961 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2960 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2959 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2958 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2957 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2956 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2955 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2954 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2953 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2952 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2951 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2950 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2949 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2948 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2947 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2946 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2945 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2944 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2943 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2942 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2941 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2940 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2939 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2938 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2937 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2936 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2935 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2934 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2933 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2932 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2931 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2930 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2929 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2928 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2927 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2926 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2925 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2924 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2923 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2922 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2921 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2920 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2919 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2918 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2917 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2916 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2915 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2914 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2913 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2912 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2911 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2910 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2909 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2908 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2907 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2906 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2905 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2904 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2903 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2902 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2901 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2900 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2899 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2898 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2897 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2896 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2895 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2894 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2893 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2892 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2891 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2890 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2889 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2888 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2887 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2886 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2885 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2884 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2883 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2882 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2881 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2880 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2879 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2878 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2877 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2876 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2875 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2874 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2873 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2872 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2871 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2870 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2869 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2868 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2867 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2866 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2865 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2864 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2863 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2862 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2861 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2860 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2859 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2858 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2857 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2856 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2855 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2854 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2853 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2852 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2851 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2850 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2849 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2848 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2847 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2846 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2845 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2844 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2843 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2842 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2841 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2840 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2839 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2838 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2837 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2836 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2835 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2834 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2833 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2832 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2831 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2830 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2829 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2828 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2827 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2826 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2825 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2824 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2823 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2822 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2821 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2820 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2819 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2818 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2817 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2816 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2815 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2814 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2813 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2812 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2811 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2810 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2809 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2808 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2807 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2806 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2805 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2804 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2803 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2802 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2801 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2800 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2799 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2798 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2797 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2796 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2795 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2794 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2793 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2792 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2791 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2790 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2789 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2788 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2787 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2786 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2785 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2784 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2783 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2782 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2781 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2780 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2779 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2778 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2777 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2776 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2775 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2774 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2773 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2772 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2771 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2770 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2769 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2768 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2767 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2766 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2765 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2764 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2763 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2762 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2761 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2760 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2759 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2758 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2757 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2756 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2755 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2754 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2753 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2752 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2751 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2750 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2749 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2748 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2747 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2746 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2745 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2744 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2743 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2742 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2741 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2740 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2739 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2738 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2737 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2736 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2735 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2734 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2733 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2732 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2731 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2730 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2729 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2728 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2727 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2726 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2725 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2724 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2723 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2722 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2721 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2720 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2719 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2718 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2717 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2716 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2715 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2714 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2713 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2712 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2711 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2710 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2709 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2708 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2707 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2706 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2705 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2704 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2703 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2702 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2701 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2700 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2699 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2698 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2697 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2696 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2695 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2694 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2693 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2692 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2691 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2690 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2689 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2688 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2687 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2686 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2685 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2684 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2683 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2682 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2681 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2680 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2679 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2678 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2677 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2676 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2675 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2674 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2673 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2672 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2671 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2670 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2669 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2668 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2667 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2666 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2665 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2664 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2663 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2662 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2661 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2660 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2659 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2658 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2657 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2656 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2655 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2654 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2653 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2652 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2651 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2650 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2649 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2648 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2647 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2646 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2645 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2644 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2643 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2642 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2641 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2640 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2639 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2638 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2637 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2636 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2635 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2634 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2633 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2632 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2631 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2630 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2629 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2628 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2627 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2626 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2625 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2624 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2623 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2622 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2621 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2620 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2619 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2618 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2617 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2616 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2615 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2614 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2613 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2612 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2611 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2610 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2609 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2608 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2607 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2606 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2605 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2604 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2603 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2602 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2601 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2600 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2599 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2598 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2597 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2596 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2595 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2594 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2593 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2592 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2591 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2590 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2589 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2588 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2587 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2586 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2585 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2584 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2583 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2582 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2581 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2580 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2579 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2578 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2577 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2576 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2575 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2574 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2573 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2572 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2571 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2570 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2569 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2568 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2567 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2566 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2565 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2564 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2563 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2562 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2561 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2560 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2559 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2558 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2557 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2556 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2555 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2554 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2553 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2552 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2551 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2550 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2549 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2548 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2547 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2546 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2545 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2544 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2543 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2542 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2541 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2540 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2539 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2538 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2537 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2536 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2535 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2534 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2533 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2532 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2531 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2530 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2529 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2528 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2527 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2526 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2525 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2524 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2523 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2522 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2521 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2520 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2519 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2518 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2517 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2516 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2515 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2514 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2513 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2512 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2511 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2510 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2509 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2508 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2507 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2506 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2505 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2504 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2503 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2502 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2501 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2500 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2499 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2498 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2497 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2496 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2495 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2494 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2493 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2492 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2491 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2490 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2489 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2488 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2487 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2486 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2485 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2484 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2483 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2482 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2481 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2480 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2479 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2478 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2477 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2476 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2475 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2474 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2473 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2472 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2471 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2470 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2469 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2468 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2467 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2466 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2465 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2464 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2463 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2462 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2461 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2460 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2459 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2458 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2457 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2456 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2455 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2454 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2453 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2452 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2451 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2450 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2449 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2448 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2447 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2446 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2445 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2444 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2443 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2442 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2441 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2440 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2439 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2438 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2437 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2436 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2435 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2434 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2433 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2432 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2431 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2430 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2429 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2428 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2427 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2426 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2425 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2424 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2423 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2422 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2421 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2420 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2419 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2418 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2417 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2416 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2415 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2414 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2413 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2412 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2411 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2410 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2409 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2408 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2407 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2406 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2405 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2404 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2403 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2402 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2401 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2400 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2399 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2398 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2397 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2396 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2395 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2394 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2393 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2392 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2391 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2390 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2389 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2388 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2387 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2386 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2385 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2384 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2383 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2382 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2381 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2380 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2379 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2378 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2377 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2376 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2375 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2374 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2373 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2372 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2371 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2370 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2369 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2368 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2367 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2366 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2365 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2364 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2363 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2362 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2361 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2360 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2359 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2358 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2357 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2356 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2355 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2354 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2353 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2352 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2351 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2350 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2349 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2348 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2347 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2346 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2345 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2344 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2343 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2342 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2341 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2340 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2339 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2338 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2337 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2336 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2335 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2334 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2333 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2332 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2331 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2330 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2329 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2328 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2327 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2326 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2325 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2324 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2323 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2322 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2321 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2320 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2319 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2318 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2317 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2316 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2315 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2314 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2313 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2312 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2311 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2310 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2309 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2308 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2307 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2306 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2305 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2304 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2303 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2302 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2301 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2300 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2299 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2298 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2297 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2296 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2295 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2294 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2293 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2292 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2291 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2290 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2289 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2288 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2287 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2286 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2285 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2284 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2283 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2282 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2281 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2280 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2279 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2278 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2277 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2276 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2275 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2274 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2273 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2272 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2271 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2270 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2269 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2268 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2267 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2266 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2265 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2264 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2263 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2262 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2261 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2260 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2259 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2258 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2257 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2256 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2255 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2254 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2253 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2252 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2251 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2250 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2249 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2248 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2247 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2246 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2245 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2244 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2243 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2242 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2241 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2240 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2239 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2238 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2237 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2236 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2235 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2234 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2233 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2232 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2231 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2230 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2229 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2228 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2227 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2226 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2225 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2224 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2223 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2222 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2221 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2220 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2219 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2218 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2217 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2216 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2215 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2214 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2213 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2212 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2211 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2210 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2209 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2208 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2207 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2206 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2205 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2204 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2203 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2202 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2201 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2200 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2199 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2198 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2197 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2196 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2195 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2194 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2193 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2192 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2191 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2190 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2189 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2188 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2187 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2186 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2185 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2184 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2183 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2182 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2181 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2180 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2179 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2178 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2177 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2176 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2175 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2174 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2173 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2172 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2171 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2170 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2169 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2168 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2167 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2166 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2165 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2164 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2163 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2162 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2161 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2160 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2159 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2158 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2157 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2156 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2155 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2154 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2153 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2152 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2151 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2150 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2149 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2148 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2147 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2146 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2145 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2144 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2143 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2142 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2141 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2140 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2139 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2138 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2137 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2136 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2135 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2134 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2133 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2132 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2131 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2130 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2129 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2128 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2127 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2126 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2125 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2124 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2123 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2122 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2121 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2120 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2119 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2118 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2117 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2116 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2115 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2114 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2113 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2112 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2111 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2110 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2109 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2108 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2107 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2106 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2105 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2104 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2103 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2102 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2101 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2100 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2099 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2098 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2097 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2096 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2095 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2094 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2093 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2092 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2091 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2090 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2089 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2088 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2087 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2086 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2085 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2084 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2083 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2082 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2081 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2080 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2079 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2078 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2077 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2076 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2075 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2074 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2073 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2072 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2071 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2070 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2069 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2068 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2067 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2066 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2065 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2064 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2063 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2062 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2061 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2060 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2059 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2058 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2057 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2056 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2055 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2054 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2053 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2052 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2051 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2050 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2049 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2048 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2047 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2046 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2045 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2044 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2043 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2042 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2041 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2040 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2039 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2038 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2037 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2036 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2035 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2034 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2033 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2032 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2031 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2030 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2029 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2028 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2027 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2026 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2025 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2024 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2023 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2022 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2021 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2020 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2019 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2018 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2017 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2016 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2015 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2014 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2013 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2012 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2011 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2010 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2009 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2008 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2007 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2006 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2005 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2004 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2003 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2002 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2001 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2000 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1999 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1998 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1997 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1996 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1995 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1994 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1993 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1992 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1991 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1990 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1989 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1988 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1987 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1986 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1985 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1984 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1983 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1982 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1981 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1980 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1979 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1978 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1977 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1976 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1975 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1974 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1973 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1972 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1971 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1970 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1969 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1968 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1967 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1966 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1965 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1964 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1963 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1962 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1961 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1960 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1959 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1958 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1957 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1956 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1955 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1954 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1953 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1952 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1951 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1950 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1949 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1948 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1947 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1946 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1945 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1944 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1943 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1942 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1941 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1940 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1939 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1938 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1937 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1936 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1935 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1934 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1933 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1932 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1931 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1930 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1929 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1928 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1927 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1926 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1925 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1924 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1923 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1922 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1921 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1920 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1919 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1918 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1917 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1916 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1915 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1914 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1913 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1912 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1911 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1910 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1909 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1908 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1907 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1906 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1905 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1904 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1903 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1902 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1901 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1900 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1899 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1898 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1897 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1896 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1895 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1894 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1893 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1892 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1891 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1890 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1889 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1888 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1887 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1886 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1885 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1884 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1883 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1882 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1881 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1880 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1879 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1878 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1877 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1876 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1875 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1874 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1873 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1872 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1871 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1870 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1869 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1868 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1867 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1866 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1865 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1864 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1863 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1862 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1861 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1860 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1859 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1858 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1857 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1856 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1855 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1854 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1853 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1852 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1851 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1850 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1849 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1848 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1847 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1846 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1845 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1844 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1843 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1842 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1841 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1840 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1839 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1838 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1837 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1836 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1835 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1834 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1833 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1832 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1831 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1830 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1829 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1828 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1827 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1826 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1825 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1824 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1823 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1822 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1821 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1820 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1819 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1818 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1817 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1816 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1815 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1814 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1813 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1812 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1811 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1810 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1809 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1808 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1807 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1806 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1805 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1804 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1803 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1802 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1801 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1800 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1799 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1798 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1797 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1796 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1795 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1794 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1793 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1792 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1791 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1790 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1789 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1788 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1787 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1786 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1785 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1784 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1783 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1782 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1781 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1780 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1779 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1778 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1777 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1776 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1775 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1774 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1773 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1772 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1771 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1770 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1769 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1768 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1767 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1766 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1765 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1764 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1763 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1762 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1761 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1760 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1759 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1758 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1757 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1756 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1755 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1754 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1753 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1752 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1751 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1750 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1749 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1748 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1747 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1746 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1745 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1744 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1743 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1742 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1741 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1740 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1739 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1738 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1737 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1736 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1735 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1734 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1733 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1732 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1731 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1730 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1729 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1728 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1727 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1726 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1725 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1724 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1723 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1722 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1721 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1720 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1719 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1718 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1717 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1716 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1715 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1714 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1713 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1712 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1711 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1710 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1709 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1708 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1707 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1706 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1705 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1704 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1703 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1702 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1701 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1700 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1699 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1698 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1697 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1696 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1695 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1694 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1693 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1692 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1691 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1690 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1689 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1688 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1687 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1686 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1685 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1684 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1683 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1682 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1681 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1680 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1679 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1678 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1677 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1676 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1675 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1674 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1673 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1672 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1671 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1670 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1669 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1668 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1667 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1666 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1665 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1664 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1663 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1662 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1661 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1660 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1659 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1658 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1657 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1656 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1655 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1654 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1653 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1652 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1651 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1650 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1649 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1648 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1647 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1646 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1645 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1644 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1643 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1642 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1641 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1640 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1639 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1638 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1637 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1636 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1635 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1634 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1633 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1632 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1631 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1630 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1629 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1628 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1627 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1626 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1625 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1624 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1623 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1622 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1621 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1620 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1619 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1618 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1617 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1616 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1615 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1614 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1613 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1612 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1611 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1610 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1609 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1608 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1607 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1606 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1605 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1604 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1603 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1602 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1601 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1600 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1599 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1598 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1597 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1596 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1595 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1594 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1593 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1592 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1591 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1590 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1589 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1588 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1587 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1586 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1585 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1584 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1583 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1582 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1581 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1580 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1579 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1578 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1577 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1576 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1575 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1574 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1573 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1572 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1571 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1570 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1569 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1568 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1567 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1566 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1565 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1564 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1563 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1562 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1561 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1560 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1559 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1558 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1557 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1556 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1555 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1554 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1553 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1552 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1551 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1550 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1549 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1548 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1547 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1546 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1545 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1544 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1543 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1542 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1541 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1540 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1539 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1538 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1537 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1536 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1535 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1534 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1533 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1532 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1531 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1530 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1529 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1528 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1527 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1526 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1525 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1524 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1523 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1522 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1521 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1520 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1519 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1518 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1517 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1516 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1515 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1514 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1513 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1512 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1511 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1510 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1509 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1508 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1507 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1506 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1505 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1504 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1503 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1502 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1501 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1500 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1499 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1498 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1497 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1496 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1495 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1494 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1493 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1492 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1491 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1490 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1489 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1488 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1487 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1486 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1485 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1484 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1483 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1482 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1481 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1480 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1479 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1478 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1477 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1476 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1475 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1474 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1473 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1472 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1471 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1470 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1469 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1468 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1467 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1466 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1465 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1464 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1463 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1462 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1461 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1460 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1459 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1458 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1457 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1456 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1455 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1454 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1453 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1452 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1451 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1450 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1449 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1448 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1447 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1446 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1445 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1444 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1443 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1442 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1441 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1440 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1439 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1438 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1437 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1436 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1435 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1434 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1433 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1432 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1431 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1430 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1429 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1428 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1427 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1426 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1425 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1424 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1423 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1422 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1421 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1420 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1419 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1418 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1417 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1416 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1415 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1414 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1413 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1412 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1411 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1410 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1409 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1408 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1407 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1406 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1405 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1404 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1403 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1402 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1401 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1400 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1399 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1398 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1397 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1396 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1395 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1394 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1393 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1392 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1391 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1390 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1389 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1388 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1387 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1386 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1385 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1384 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1383 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1382 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1381 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1380 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1379 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1378 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1377 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1376 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1375 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1374 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1373 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1372 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1371 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1370 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1369 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1368 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1367 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1366 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1365 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1364 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1363 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1362 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1361 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1360 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1359 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1358 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1357 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1356 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1355 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1354 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1353 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1352 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1351 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1350 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1349 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1348 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1347 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1346 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1345 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1344 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1343 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1342 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1341 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1340 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1339 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1338 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1337 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1336 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1335 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1334 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1333 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1332 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1331 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1330 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1329 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1328 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1327 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1326 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1325 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1324 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1323 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1322 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1321 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1320 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1319 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1318 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1317 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1316 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1315 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1314 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1313 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1312 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1311 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1310 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1309 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1308 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1307 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1306 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1305 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1304 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1303 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1302 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1301 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1300 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1299 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1298 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1297 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1296 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1295 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1294 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1293 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1292 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1291 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1290 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1289 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1288 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1287 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1286 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1285 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1284 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1283 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1282 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1281 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1280 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1279 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1278 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1277 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1276 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1275 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1274 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1273 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1272 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1271 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1270 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1269 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1268 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1267 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1266 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1265 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1264 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1263 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1262 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1261 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1260 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1259 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1258 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1257 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1256 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1255 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1254 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1253 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1252 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1251 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1250 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1249 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1248 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1247 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1246 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1245 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1244 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1243 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1242 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1241 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1240 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1239 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1238 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1237 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1236 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1235 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1234 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1233 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1232 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1231 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1230 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1229 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1228 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1227 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1226 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1225 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1224 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1223 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1222 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1221 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1220 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1219 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1218 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1217 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1216 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1215 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1214 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1213 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1212 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1211 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1210 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1209 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1208 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1207 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1206 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1205 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1204 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1203 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1202 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1201 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1200 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1199 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1198 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1197 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1196 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1195 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1194 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1193 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1192 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1191 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1190 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1189 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1188 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1187 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1186 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1185 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1184 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1183 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1182 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1181 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1180 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1179 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1178 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1177 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1176 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1175 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1174 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1173 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1172 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1171 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1170 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1169 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1168 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1167 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1166 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1165 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1164 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1163 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1162 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1161 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1160 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1159 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1158 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1157 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1156 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1155 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1154 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1153 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1152 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1151 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1150 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1149 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1148 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1147 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1146 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1145 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1144 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1143 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1142 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1141 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1140 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1139 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1138 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1137 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1136 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1135 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1134 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1133 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1132 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1131 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1130 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1129 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1128 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1127 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1126 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1125 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1124 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1123 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1122 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1121 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1120 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1119 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1118 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1117 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1116 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1115 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1114 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1113 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1112 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1111 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1110 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1109 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1108 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1107 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1106 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1105 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1104 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1103 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1102 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1101 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1100 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1099 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1098 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1097 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1096 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1095 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1094 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1093 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1092 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1091 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1090 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1089 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1088 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1087 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1086 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1085 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1084 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1083 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1082 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1081 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1080 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1079 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1078 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1077 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1076 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1075 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1074 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1073 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1072 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1071 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1070 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1069 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1068 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1067 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1066 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1065 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1064 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1063 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1062 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1061 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1060 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1059 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1058 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1057 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1056 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1055 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1054 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1053 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1052 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1051 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1050 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1049 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1048 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1047 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1046 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1045 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1044 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1043 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1042 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1041 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1040 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1039 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1038 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1037 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1036 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1035 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1034 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1033 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1032 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1031 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1030 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1029 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1028 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1027 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1026 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1025 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1024 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1023 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1022 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1021 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1020 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1019 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1018 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1017 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1016 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1015 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1014 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1013 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1012 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1011 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1010 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1009 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1008 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1007 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1006 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1005 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1004 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1003 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1002 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1001 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1000 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_999 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_998 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_997 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_996 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_995 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_994 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_993 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_992 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_991 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_990 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_989 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_988 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_987 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_986 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_985 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_984 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_983 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_982 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_981 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_980 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_979 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_978 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_977 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_976 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_975 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_974 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_973 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_972 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_971 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_970 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_969 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_968 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_967 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_966 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_965 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_964 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_963 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_962 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_961 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_960 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_959 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_958 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_957 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_956 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_955 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_954 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_953 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_952 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_951 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_950 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_949 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_948 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_947 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_946 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_945 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_944 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_943 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_942 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_941 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_940 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_939 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_938 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_937 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_936 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_935 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_934 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_933 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_932 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_931 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_930 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_929 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_928 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_927 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_926 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_925 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_924 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_923 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_922 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_921 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_920 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_919 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_918 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_917 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_916 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_915 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_914 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_913 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_912 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_911 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_910 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_909 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_908 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_907 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_906 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_905 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_904 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_903 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_902 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_901 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_900 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_899 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_898 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_897 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_896 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_895 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_894 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_893 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_892 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_891 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_890 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_889 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_888 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_887 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_886 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_885 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_884 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_883 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_882 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_881 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_880 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_879 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_878 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_877 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_876 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_875 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_874 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_873 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_872 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_871 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_870 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_869 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_868 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_867 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_866 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_865 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_864 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_863 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_862 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_861 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_860 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_859 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_858 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_857 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_856 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_855 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_854 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_853 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_852 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_851 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_850 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_849 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_848 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_847 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_846 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_845 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_844 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_843 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_842 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_841 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_840 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_839 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_838 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_837 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_836 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_835 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_834 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_833 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_832 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_831 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_830 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_829 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_828 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_827 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_826 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_825 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_824 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_823 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_822 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_821 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_820 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_819 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_818 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_817 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_816 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_815 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_814 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_813 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_812 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_811 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_810 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_809 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_808 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_807 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_806 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_805 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_804 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_803 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_802 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_801 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_800 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_799 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_798 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_797 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_796 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_795 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_794 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_793 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_792 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_791 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_790 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_789 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_788 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_787 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_786 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_785 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_784 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_783 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_782 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_781 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_780 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_779 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_778 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_777 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_776 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_775 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_774 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_773 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_772 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_771 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_770 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_769 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_768 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_767 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_766 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_765 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_764 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_763 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_762 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_761 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_760 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_759 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_758 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_757 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_756 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_755 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_754 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_753 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_752 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_751 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_750 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_749 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_748 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_747 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_746 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_745 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_744 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_743 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_742 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_741 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_740 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_739 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_738 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_737 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_736 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_735 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_734 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_733 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_732 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_731 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_730 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_729 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_728 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_727 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_726 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_725 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_724 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_723 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_722 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_721 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_720 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_719 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_718 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_717 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_716 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_715 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_714 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_713 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_712 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_711 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_710 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_709 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_708 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_707 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_706 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_705 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_704 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_703 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_702 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_701 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_700 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_699 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_698 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_697 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_696 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_695 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_694 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_693 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_692 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_691 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_690 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_689 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_688 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_687 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_686 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_685 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_684 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_683 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_682 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_681 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_680 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_679 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_678 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_677 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_676 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_675 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_674 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_673 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_672 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_671 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_670 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_669 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_668 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_667 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_666 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X4 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(N1) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X4 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X4 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X2 U1 ( .A(A), .ZN(Y) );
endmodule


module Sum_generator_Nbit32_Nblock8_6 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_48 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  cs_generic_N4_47 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  cs_generic_N4_46 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  cs_generic_N4_45 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_44 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_43 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_42 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_41 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module Sum_generator_Nbit32_Nblock8_5 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_40 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  cs_generic_N4_39 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  cs_generic_N4_38 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  cs_generic_N4_37 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_36 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_35 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_34 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_33 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module Sum_generator_Nbit32_Nblock8_4 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_32 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  cs_generic_N4_31 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  cs_generic_N4_30 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  cs_generic_N4_29 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_28 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_27 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_26 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_25 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module Sum_generator_Nbit32_Nblock8_3 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_24 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  cs_generic_N4_23 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  cs_generic_N4_22 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  cs_generic_N4_21 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_20 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_19 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_18 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_17 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module Sum_generator_Nbit32_Nblock8_2 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_16 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0])
         );
  cs_generic_N4_15 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  cs_generic_N4_14 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  cs_generic_N4_13 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_12 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_11 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_10 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_9 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module Sum_generator_Nbit32_Nblock8_1 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_8 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  cs_generic_N4_7 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  cs_generic_N4_6 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  cs_generic_N4_5 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_4 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_3 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_2 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_1 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sparce_tree_POWER5_6 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] , n1, n2, n3,
         n4, n5, n6;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U46 ( .A(B[28]), .B(A[28]), .Z(\matrixP[28][28] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_60 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_59 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_162 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), 
        .Gik(\matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), 
        .Gij(\matrixG[4][3] ) );
  block_pg_161 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), 
        .Gik(\matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), 
        .Gij(\matrixG[6][5] ) );
  block_pg_160 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), 
        .Gik(\matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), 
        .Gij(\matrixG[8][7] ) );
  block_pg_159 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_158 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_157 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_156 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_155 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_154 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_153 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_152 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_151 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_150 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_149 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_148 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_58 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_147 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), 
        .Gik(\matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), 
        .Gij(\matrixG[8][5] ) );
  block_pg_146 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_145 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_144 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_143 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_142 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_141 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_57 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_140 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_139 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(n2), .Pij(\matrixP[24][17] ), .Gij(
        \matrixG[24][17] ) );
  block_pg_138 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_56 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_55 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_137 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_136 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_54 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_53 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_52 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_51 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  NAND2_X2 U1 ( .A1(n4), .A2(n5), .ZN(\matrixP[20][20] ) );
  INV_X2 U2 ( .A(B[20]), .ZN(n3) );
  INV_X1 U3 ( .A(A[16]), .ZN(n1) );
  AND2_X2 U4 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  XOR2_X2 U5 ( .A(B[24]), .B(A[24]), .Z(\matrixP[24][24] ) );
  XNOR2_X2 U6 ( .A(B[16]), .B(n1), .ZN(\matrixP[16][16] ) );
  NAND2_X1 U7 ( .A1(n3), .A2(A[20]), .ZN(n5) );
  AND2_X1 U8 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U9 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  AND2_X1 U10 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U11 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U12 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U13 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U14 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  INV_X1 U15 ( .A(A[20]), .ZN(n6) );
  AND2_X1 U16 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U17 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  AND2_X1 U18 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U19 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U20 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U21 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U22 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U23 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U24 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U25 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U26 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
  AND2_X1 U27 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U28 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U29 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U30 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U31 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U32 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U50 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U54 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U58 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U65 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U66 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  AND2_X1 U67 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  CLKBUF_X1 U68 ( .A(\matrixG[20][17] ), .Z(n2) );
  NAND2_X1 U69 ( .A1(B[20]), .A2(n6), .ZN(n4) );
  AND2_X1 U70 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
endmodule


module sparce_tree_POWER5_5 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] , n1, n2, n3,
         n4;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U46 ( .A(B[28]), .B(A[28]), .Z(\matrixP[28][28] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_50 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_49 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_135 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), 
        .Gik(\matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), 
        .Gij(\matrixG[4][3] ) );
  block_pg_134 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), 
        .Gik(\matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), 
        .Gij(\matrixG[6][5] ) );
  block_pg_133 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), 
        .Gik(\matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), 
        .Gij(\matrixG[8][7] ) );
  block_pg_132 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_131 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_130 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_129 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_128 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_127 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_126 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_125 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_124 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_123 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_122 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_121 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_48 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_120 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), 
        .Gik(\matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), 
        .Gij(\matrixG[8][5] ) );
  block_pg_119 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_118 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_117 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_116 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_115 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_114 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_47 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_113 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_112 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_111 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_46 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_45 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_110 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_109 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_44 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_43 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_42 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_41 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(\matrixP[20][20] ) );
  NAND2_X1 U2 ( .A1(B[20]), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A[20]), .ZN(n4) );
  INV_X1 U4 ( .A(B[20]), .ZN(n1) );
  INV_X1 U5 ( .A(A[20]), .ZN(n2) );
  XOR2_X1 U6 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U7 ( .A(B[24]), .B(A[24]), .Z(\matrixP[24][24] ) );
  XOR2_X1 U8 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  AND2_X1 U9 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
  AND2_X1 U10 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U11 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U12 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  AND2_X1 U13 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U14 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U15 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  AND2_X1 U16 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  AND2_X1 U17 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U18 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U19 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U20 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U21 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U22 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U23 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U24 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U25 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U26 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U27 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U28 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
  AND2_X1 U29 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U31 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U32 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U50 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U54 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U58 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U62 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U65 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U66 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  AND2_X1 U67 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  AND2_X1 U68 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
endmodule


module sparce_tree_POWER5_4 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] , n1, n2, n3,
         n4, n5, n6, n7, n8;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_40 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_39 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_108 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), 
        .Gik(\matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), 
        .Gij(\matrixG[4][3] ) );
  block_pg_107 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), 
        .Gik(\matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), 
        .Gij(\matrixG[6][5] ) );
  block_pg_106 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), 
        .Gik(\matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), 
        .Gij(\matrixG[8][7] ) );
  block_pg_105 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_104 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_103 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_102 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_101 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_100 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_99 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_98 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_97 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_96 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_95 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_94 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_38 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_93 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), .Gik(
        \matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), .Gij(
        \matrixG[8][5] ) );
  block_pg_92 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_91 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_90 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_89 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_88 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_87 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_37 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_86 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_85 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_84 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_36 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_35 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_83 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_82 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_34 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_33 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_32 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_31 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  XOR2_X2 U1 ( .A(B[28]), .B(A[28]), .Z(\matrixP[28][28] ) );
  AND2_X2 U2 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  NAND2_X1 U3 ( .A1(B[24]), .A2(n8), .ZN(n6) );
  INV_X1 U4 ( .A(B[20]), .ZN(n1) );
  NAND2_X2 U5 ( .A1(n5), .A2(A[24]), .ZN(n7) );
  NAND2_X2 U6 ( .A1(n6), .A2(n7), .ZN(\matrixP[24][24] ) );
  AND2_X2 U7 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  NAND2_X1 U8 ( .A1(n2), .A2(n3), .ZN(\matrixP[20][20] ) );
  NAND2_X1 U9 ( .A1(n1), .A2(A[20]), .ZN(n3) );
  XOR2_X1 U10 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  AND2_X1 U11 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U12 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U13 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U14 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U15 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  INV_X1 U16 ( .A(A[20]), .ZN(n4) );
  INV_X1 U17 ( .A(A[24]), .ZN(n8) );
  AND2_X1 U18 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U19 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U20 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U21 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U22 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U23 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U24 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U25 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U26 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U27 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U28 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U29 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
  AND2_X1 U30 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U31 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U32 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U46 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U50 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U54 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U58 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U65 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U66 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U67 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  NAND2_X1 U68 ( .A1(B[20]), .A2(n4), .ZN(n2) );
  AND2_X1 U69 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  INV_X1 U70 ( .A(B[24]), .ZN(n5) );
  AND2_X1 U71 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
  AND2_X1 U72 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
endmodule


module sparce_tree_POWER5_3 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] , n1;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_30 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_29 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_81 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), .Gik(
        \matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), .Gij(
        \matrixG[4][3] ) );
  block_pg_80 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), .Gik(
        \matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), .Gij(
        \matrixG[6][5] ) );
  block_pg_79 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), .Gik(
        \matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), .Gij(
        \matrixG[8][7] ) );
  block_pg_78 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_77 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_76 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_75 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_74 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_73 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_72 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_71 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_70 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_69 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_68 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_67 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_28 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_66 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), .Gik(
        \matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), .Gij(
        \matrixG[8][5] ) );
  block_pg_65 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_64 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_63 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_62 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_61 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_60 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_27 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_59 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_58 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_57 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_26 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_25 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_56 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_55 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_24 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_23 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_22 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_21 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  INV_X1 U1 ( .A(A[24]), .ZN(n1) );
  XOR2_X2 U2 ( .A(B[28]), .B(A[28]), .Z(\matrixP[28][28] ) );
  XNOR2_X2 U3 ( .A(B[24]), .B(n1), .ZN(\matrixP[24][24] ) );
  XOR2_X1 U4 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  XOR2_X1 U5 ( .A(B[20]), .B(A[20]), .Z(\matrixP[20][20] ) );
  AND2_X1 U6 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U7 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U8 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U9 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U10 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  AND2_X1 U11 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U12 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  AND2_X1 U13 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U14 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  AND2_X1 U15 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U16 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U17 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U18 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  AND2_X1 U19 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U20 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U21 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U22 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U23 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U24 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U25 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U26 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U27 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U28 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U29 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U30 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U31 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U32 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U46 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U50 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
  AND2_X1 U54 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  AND2_X1 U58 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  AND2_X1 U65 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
endmodule


module sparce_tree_POWER5_2 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] , n1, n2, n3,
         n4, n5;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U54 ( .A(B[20]), .B(A[20]), .Z(\matrixP[20][20] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U58 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_20 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_19 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_54 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), .Gik(
        \matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), .Gij(
        \matrixG[4][3] ) );
  block_pg_53 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), .Gik(
        \matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), .Gij(
        \matrixG[6][5] ) );
  block_pg_52 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), .Gik(
        \matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), .Gij(
        \matrixG[8][7] ) );
  block_pg_51 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_50 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_49 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_48 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_47 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_46 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_45 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_44 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_43 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_42 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_41 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_40 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_18 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_39 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), .Gik(
        \matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), .Gij(
        \matrixG[8][5] ) );
  block_pg_38 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_37 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_36 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_35 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_34 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_33 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_17 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_32 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_31 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_30 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_16 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_15 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_29 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_28 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_14 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_13 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_12 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_11 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  XNOR2_X2 U1 ( .A(B[28]), .B(n1), .ZN(\matrixP[28][28] ) );
  INV_X1 U2 ( .A(A[28]), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n4), .A2(n5), .ZN(\matrixP[24][24] ) );
  NAND2_X1 U4 ( .A1(B[24]), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n2), .A2(A[24]), .ZN(n5) );
  INV_X1 U6 ( .A(B[24]), .ZN(n2) );
  INV_X1 U7 ( .A(A[24]), .ZN(n3) );
  XOR2_X1 U8 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  AND2_X1 U9 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U10 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U11 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U12 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U13 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  AND2_X1 U14 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  AND2_X1 U15 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  AND2_X1 U16 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  AND2_X1 U17 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U18 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  AND2_X1 U19 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U20 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U21 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U22 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
  AND2_X1 U23 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U24 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U25 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U26 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U27 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U28 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U29 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U30 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U31 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U32 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U46 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U48 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U50 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U65 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  AND2_X1 U66 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U67 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U68 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U69 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
endmodule


module sparce_tree_POWER5_1 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] , n1;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U54 ( .A(B[20]), .B(A[20]), .Z(\matrixP[20][20] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U58 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_10 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_9 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_27 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), .Gik(
        \matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), .Gij(
        \matrixG[4][3] ) );
  block_pg_26 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), .Gik(
        \matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), .Gij(
        \matrixG[6][5] ) );
  block_pg_25 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), .Gik(
        \matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), .Gij(
        \matrixG[8][7] ) );
  block_pg_24 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_23 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_22 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_21 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_20 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_19 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_18 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_17 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_16 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_15 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_14 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_13 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_8 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_12 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), .Gik(
        \matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), .Gij(
        \matrixG[8][5] ) );
  block_pg_11 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_10 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_9 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_8 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_7 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_6 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_7 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_5 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_4 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_3 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_6 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_5 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_2 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_1 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_4 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_3 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_2 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_1 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  XNOR2_X1 U1 ( .A(B[28]), .B(n1), .ZN(\matrixP[28][28] ) );
  INV_X1 U2 ( .A(A[28]), .ZN(n1) );
  AND2_X2 U3 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  XOR2_X1 U4 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U5 ( .A(B[24]), .B(A[24]), .Z(\matrixP[24][24] ) );
  AND2_X1 U6 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U7 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U8 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  AND2_X1 U9 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  AND2_X1 U10 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U11 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U12 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U13 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U14 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U15 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  AND2_X1 U16 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U17 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  AND2_X1 U18 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U19 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U20 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U21 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U22 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U23 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
  AND2_X1 U24 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U25 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
  AND2_X1 U26 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U28 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U30 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  AND2_X1 U31 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U32 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U46 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U50 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U52 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U65 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
endmodule


module MUX21_GENERIC_N32_31 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_87 UIV ( .A(n1), .Y(SB) );
  ND2_3648 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3647 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_3646 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3645 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3644 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_3643 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3642 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3641 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_3640 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3639 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3638 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_3637 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3636 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3635 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_3634 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3633 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3632 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_3631 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3630 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3629 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_3628 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3627 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3626 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_3625 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3624 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3623 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_3622 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3621 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3620 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_3619 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3618 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3617 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_3616 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3615 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3614 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_3613 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3612 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3611 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_3610 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3609 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3608 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_3607 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3606 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3605 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_3604 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3603 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3602 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_3601 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3600 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3599 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_3598 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3597 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3596 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_3595 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3594 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3593 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_3592 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3591 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3590 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3589 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3588 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3587 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3586 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3585 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3584 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3583 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3582 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3581 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3580 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3579 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3578 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_3577 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3576 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3575 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_3574 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3573 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3572 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_3571 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3570 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3569 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_3568 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3567 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3566 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_3565 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3564 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3563 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_3562 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3561 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3560 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_3559 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3558 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3557 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_3556 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3555 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3554 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_3553 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  CLKBUF_X1 U1 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U2 ( .A(SEL), .Z(n3) );
  CLKBUF_X1 U3 ( .A(SB), .Z(n5) );
  CLKBUF_X1 U4 ( .A(SB), .Z(n6) );
  BUF_X1 U5 ( .A(SB), .Z(n4) );
  BUF_X2 U6 ( .A(SEL), .Z(n1) );
endmodule


module MUX21_GENERIC_N32_30 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_86 UIV ( .A(n1), .Y(SB) );
  ND2_3552 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3551 UND2_31 ( .A(B[31]), .B(n5), .Y(Y2[31]) );
  ND2_3550 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3549 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3548 UND2_30 ( .A(B[30]), .B(n5), .Y(Y2[30]) );
  ND2_3547 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3546 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3545 UND2_29 ( .A(B[29]), .B(n5), .Y(Y2[29]) );
  ND2_3544 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3543 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3542 UND2_28 ( .A(B[28]), .B(n5), .Y(Y2[28]) );
  ND2_3541 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3540 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3539 UND2_27 ( .A(B[27]), .B(n5), .Y(Y2[27]) );
  ND2_3538 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3537 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3536 UND2_26 ( .A(B[26]), .B(n5), .Y(Y2[26]) );
  ND2_3535 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3534 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3533 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  ND2_3532 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3531 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3530 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  ND2_3529 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3528 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3527 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  ND2_3526 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3525 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3524 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  ND2_3523 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3522 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3521 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  ND2_3520 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3519 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3518 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  ND2_3517 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3516 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3515 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  ND2_3514 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3513 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3512 UND2_18 ( .A(B[18]), .B(n4), .Y(Y2[18]) );
  ND2_3511 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3510 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3509 UND2_17 ( .A(B[17]), .B(n4), .Y(Y2[17]) );
  ND2_3508 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3507 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3506 UND2_16 ( .A(B[16]), .B(n4), .Y(Y2[16]) );
  ND2_3505 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3504 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3503 UND2_15 ( .A(B[15]), .B(n4), .Y(Y2[15]) );
  ND2_3502 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3501 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3500 UND2_14 ( .A(B[14]), .B(n4), .Y(Y2[14]) );
  ND2_3499 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3498 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3497 UND2_13 ( .A(B[13]), .B(n4), .Y(Y2[13]) );
  ND2_3496 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3495 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3494 UND2_12 ( .A(B[12]), .B(SB), .Y(Y2[12]) );
  ND2_3493 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3492 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3491 UND2_11 ( .A(B[11]), .B(SB), .Y(Y2[11]) );
  ND2_3490 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3489 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3488 UND2_10 ( .A(B[10]), .B(SB), .Y(Y2[10]) );
  ND2_3487 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3486 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3485 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3484 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3483 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3482 UND2_8 ( .A(B[8]), .B(SB), .Y(Y2[8]) );
  ND2_3481 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3480 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3479 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  ND2_3478 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3477 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3476 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_3475 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3474 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3473 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  ND2_3472 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3471 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3470 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  ND2_3469 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3468 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3467 UND2_3 ( .A(B[3]), .B(n5), .Y(Y2[3]) );
  ND2_3466 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3465 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3464 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_3463 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3462 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3461 UND2_1 ( .A(B[1]), .B(n5), .Y(Y2[1]) );
  ND2_3460 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3459 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3458 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_3457 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X2 U3 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U4 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U5 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_29 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_85 UIV ( .A(n1), .Y(SB) );
  ND2_3456 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3455 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_3454 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3453 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3452 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_3451 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3450 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3449 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_3448 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3447 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3446 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_3445 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3444 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3443 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_3442 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3441 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3440 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_3439 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3438 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3437 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_3436 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3435 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3434 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_3433 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3432 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3431 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_3430 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3429 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3428 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_3427 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3426 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3425 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_3424 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3423 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3422 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_3421 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3420 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3419 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_3418 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3417 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3416 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_3415 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3414 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3413 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_3412 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3411 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3410 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_3409 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3408 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3407 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_3406 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3405 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3404 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_3403 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3402 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3401 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_3400 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3399 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3398 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3397 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3396 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3395 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3394 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3393 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3392 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3391 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3390 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3389 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3388 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3387 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3386 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_3385 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3384 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3383 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_3382 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3381 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3380 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_3379 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3378 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3377 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_3376 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3375 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3374 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_3373 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3372 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3371 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_3370 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3369 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3368 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_3367 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3366 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3365 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_3364 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3363 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3362 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_3361 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U2 ( .A(SB), .Z(n5) );
  CLKBUF_X1 U3 ( .A(SB), .Z(n6) );
  CLKBUF_X1 U4 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U5 ( .A(SEL), .Z(n3) );
  BUF_X1 U6 ( .A(SB), .Z(n4) );
endmodule


module MUX21_GENERIC_N32_28 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_84 UIV ( .A(n1), .Y(SB) );
  ND2_3360 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3359 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_3358 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3357 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3356 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_3355 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3354 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3353 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_3352 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3351 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3350 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_3349 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3348 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3347 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_3346 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3345 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3344 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_3343 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3342 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3341 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_3340 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3339 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3338 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_3337 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3336 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3335 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_3334 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3333 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3332 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_3331 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3330 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3329 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_3328 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3327 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3326 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_3325 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3324 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3323 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_3322 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3321 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3320 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_3319 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3318 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3317 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_3316 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3315 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3314 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_3313 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3312 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3311 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_3310 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3309 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3308 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_3307 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3306 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3305 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_3304 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3303 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3302 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3301 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3300 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3299 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3298 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3297 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3296 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3295 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3294 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3293 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3292 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3291 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3290 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_3289 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3288 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3287 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_3286 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3285 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3284 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_3283 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3282 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3281 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_3280 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3279 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3278 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_3277 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3276 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3275 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_3274 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3273 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3272 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_3271 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3270 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3269 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_3268 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3267 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3266 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_3265 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  CLKBUF_X2 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  CLKBUF_X1 U3 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U4 ( .A(SEL), .Z(n3) );
  BUF_X1 U5 ( .A(SB), .Z(n5) );
  BUF_X1 U6 ( .A(SB), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_27 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_83 UIV ( .A(n1), .Y(SB) );
  ND2_3264 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3263 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_3262 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3261 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3260 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_3259 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3258 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3257 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_3256 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3255 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3254 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_3253 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3252 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3251 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_3250 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3249 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3248 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_3247 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3246 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3245 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_3244 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3243 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3242 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_3241 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3240 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3239 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_3238 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3237 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3236 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_3235 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3234 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3233 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_3232 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3231 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3230 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_3229 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3228 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3227 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_3226 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3225 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3224 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_3223 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3222 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3221 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_3220 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3219 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3218 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_3217 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3216 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3215 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_3214 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3213 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3212 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_3211 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3210 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3209 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_3208 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3207 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3206 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3205 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3204 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3203 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3202 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3201 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3200 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3199 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3198 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3197 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3196 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3195 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3194 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_3193 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3192 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3191 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_3190 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3189 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3188 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_3187 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3186 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3185 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_3184 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3183 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3182 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_3181 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3180 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3179 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_3178 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3177 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3176 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_3175 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3174 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3173 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_3172 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3171 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3170 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_3169 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X4 U1 ( .A(SB), .Z(n4) );
  CLKBUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X2 U3 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U4 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U5 ( .A(SEL), .Z(n3) );
  BUF_X1 U6 ( .A(SB), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_26 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_82 UIV ( .A(n1), .Y(SB) );
  ND2_3168 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3167 UND2_31 ( .A(B[31]), .B(n5), .Y(Y2[31]) );
  ND2_3166 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3165 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3164 UND2_30 ( .A(B[30]), .B(n5), .Y(Y2[30]) );
  ND2_3163 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3162 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3161 UND2_29 ( .A(B[29]), .B(n5), .Y(Y2[29]) );
  ND2_3160 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3159 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3158 UND2_28 ( .A(B[28]), .B(n5), .Y(Y2[28]) );
  ND2_3157 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3156 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3155 UND2_27 ( .A(B[27]), .B(n5), .Y(Y2[27]) );
  ND2_3154 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3153 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3152 UND2_26 ( .A(B[26]), .B(n5), .Y(Y2[26]) );
  ND2_3151 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3150 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3149 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  ND2_3148 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3147 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3146 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  ND2_3145 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3144 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3143 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  ND2_3142 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3141 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3140 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  ND2_3139 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3138 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3137 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  ND2_3136 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3135 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3134 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  ND2_3133 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3132 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3131 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  ND2_3130 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3129 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3128 UND2_18 ( .A(B[18]), .B(n4), .Y(Y2[18]) );
  ND2_3127 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3126 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3125 UND2_17 ( .A(B[17]), .B(n4), .Y(Y2[17]) );
  ND2_3124 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3123 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3122 UND2_16 ( .A(B[16]), .B(n4), .Y(Y2[16]) );
  ND2_3121 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3120 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3119 UND2_15 ( .A(B[15]), .B(n4), .Y(Y2[15]) );
  ND2_3118 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3117 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3116 UND2_14 ( .A(B[14]), .B(n4), .Y(Y2[14]) );
  ND2_3115 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3114 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3113 UND2_13 ( .A(B[13]), .B(n4), .Y(Y2[13]) );
  ND2_3112 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3111 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3110 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3109 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3108 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3107 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3106 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3105 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3104 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3103 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3102 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3101 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3100 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3099 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3098 UND2_8 ( .A(B[8]), .B(SB), .Y(Y2[8]) );
  ND2_3097 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3096 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3095 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  ND2_3094 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3093 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3092 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  ND2_3091 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3090 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3089 UND2_5 ( .A(B[5]), .B(n5), .Y(Y2[5]) );
  ND2_3088 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3087 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3086 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  ND2_3085 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3084 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3083 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_3082 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3081 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3080 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_3079 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3078 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3077 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_3076 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3075 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3074 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_3073 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X2 U2 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U3 ( .A(SB), .Z(n4) );
  CLKBUF_X1 U4 ( .A(SEL), .Z(n2) );
  CLKBUF_X1 U5 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_25 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_81 UIV ( .A(n1), .Y(SB) );
  ND2_3072 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_3071 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_3070 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3069 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3068 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_3067 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3066 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3065 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_3064 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3063 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3062 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_3061 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3060 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3059 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_3058 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3057 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3056 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_3055 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3054 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3053 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_3052 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3051 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_3050 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_3049 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3048 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3047 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_3046 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3045 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3044 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_3043 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3042 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3041 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_3040 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3039 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3038 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_3037 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3036 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3035 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_3034 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3033 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3032 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_3031 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3030 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3029 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_3028 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3027 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3026 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_3025 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3024 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3023 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_3022 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3021 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3020 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_3019 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3018 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3017 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_3016 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3015 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3014 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3013 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3012 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_3011 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3010 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3009 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3008 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3007 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3006 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3005 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3004 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3003 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3002 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_3001 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3000 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2999 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2998 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2997 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2996 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2995 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2994 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2993 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2992 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2991 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2990 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2989 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2988 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2987 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2986 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2985 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2984 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2983 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2982 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2981 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2980 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2979 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2978 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2977 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n4) );
  BUF_X1 U4 ( .A(SB), .Z(n6) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_24 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_80 UIV ( .A(n1), .Y(SB) );
  ND2_2976 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2975 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2974 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2973 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2972 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2971 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2970 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2969 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2968 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2967 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2966 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2965 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2964 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2963 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2962 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2961 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2960 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2959 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2958 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2957 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2956 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2955 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2954 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2953 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2952 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2951 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2950 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2949 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2948 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2947 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2946 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2945 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2944 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2943 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2942 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2941 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2940 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2939 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2938 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2937 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2936 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2935 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2934 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2933 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2932 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2931 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2930 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2929 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2928 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2927 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2926 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2925 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2924 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2923 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2922 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2921 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2920 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2919 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2918 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2917 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2916 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2915 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2914 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2913 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2912 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2911 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2910 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2909 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2908 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2907 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2906 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2905 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2904 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2903 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2902 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2901 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2900 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2899 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2898 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2897 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2896 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2895 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2894 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2893 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2892 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2891 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2890 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2889 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2888 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2887 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2886 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2885 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2884 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2883 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2882 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2881 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_23 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_79 UIV ( .A(n1), .Y(SB) );
  ND2_2880 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2879 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2878 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2877 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2876 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2875 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2874 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2873 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2872 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2871 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2870 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2869 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2868 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2867 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2866 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2865 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2864 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2863 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2862 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2861 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2860 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2859 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2858 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2857 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2856 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2855 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2854 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2853 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2852 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2851 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2850 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2849 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2848 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2847 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2846 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2845 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2844 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2843 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2842 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2841 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2840 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2839 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2838 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2837 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2836 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2835 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2834 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2833 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2832 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2831 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2830 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2829 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2828 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2827 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2826 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2825 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2824 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2823 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2822 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2821 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2820 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2819 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2818 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2817 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2816 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2815 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2814 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2813 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2812 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2811 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2810 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2809 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2808 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2807 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2806 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2805 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2804 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2803 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2802 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2801 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2800 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2799 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2798 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2797 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2796 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2795 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2794 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2793 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2792 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2791 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2790 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2789 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2788 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2787 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2786 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2785 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_22 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_78 UIV ( .A(n1), .Y(SB) );
  ND2_2784 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2783 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2782 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2781 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2780 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2779 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2778 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2777 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2776 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2775 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2774 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2773 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2772 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2771 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2770 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2769 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2768 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2767 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2766 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2765 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2764 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2763 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2762 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2761 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2760 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2759 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2758 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2757 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2756 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2755 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2754 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2753 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2752 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2751 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2750 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2749 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2748 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2747 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2746 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2745 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2744 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2743 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2742 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2741 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2740 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2739 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2738 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2737 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2736 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2735 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2734 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2733 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2732 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2731 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2730 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2729 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2728 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2727 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2726 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2725 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2724 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2723 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2722 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2721 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2720 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2719 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2718 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2717 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2716 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2715 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2714 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2713 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2712 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2711 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2710 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2709 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2708 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2707 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2706 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2705 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2704 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2703 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2702 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2701 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2700 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2699 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2698 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2697 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2696 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2695 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2694 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2693 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2692 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2691 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2690 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2689 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_21 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_77 UIV ( .A(n1), .Y(SB) );
  ND2_2688 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2687 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2686 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2685 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2684 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2683 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2682 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2681 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2680 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2679 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2678 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2677 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2676 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2675 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2674 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2673 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2672 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2671 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2670 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2669 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2668 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2667 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2666 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2665 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2664 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2663 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2662 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2661 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2660 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2659 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2658 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2657 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2656 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2655 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2654 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2653 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2652 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2651 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2650 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2649 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2648 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2647 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2646 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2645 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2644 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2643 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2642 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2641 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2640 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2639 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2638 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2637 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2636 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2635 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2634 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2633 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2632 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2631 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2630 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2629 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2628 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2627 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2626 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2625 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2624 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2623 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2622 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2621 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2620 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2619 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2618 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2617 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2616 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2615 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2614 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2613 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2612 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2611 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2610 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2609 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2608 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2607 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2606 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2605 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2604 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2603 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2602 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2601 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2600 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2599 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2598 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2597 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2596 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2595 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2594 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2593 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_20 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_76 UIV ( .A(n1), .Y(SB) );
  ND2_2592 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2591 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2590 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2589 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2588 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2587 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2586 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2585 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2584 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2583 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2582 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2581 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2580 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2579 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2578 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2577 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2576 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2575 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2574 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2573 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2572 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2571 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2570 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2569 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2568 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2567 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2566 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2565 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2564 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2563 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2562 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2561 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2560 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2559 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2558 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2557 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2556 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2555 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2554 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2553 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2552 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2551 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2550 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2549 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2548 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2547 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2546 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2545 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2544 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2543 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2542 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2541 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2540 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2539 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2538 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2537 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2536 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2535 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2534 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2533 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2532 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2531 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2530 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2529 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2528 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2527 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2526 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2525 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2524 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2523 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2522 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2521 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2520 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2519 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2518 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2517 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2516 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2515 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2514 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2513 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2512 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2511 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2510 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2509 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2508 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2507 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2506 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2505 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2504 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2503 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2502 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2501 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2500 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2499 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2498 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2497 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_19 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_75 UIV ( .A(n1), .Y(SB) );
  ND2_2496 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2495 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2494 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2493 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2492 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2491 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2490 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2489 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2488 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2487 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2486 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2485 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2484 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2483 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2482 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2481 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2480 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2479 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2478 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2477 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2476 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2475 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2474 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2473 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2472 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2471 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2470 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2469 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2468 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2467 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2466 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2465 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2464 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2463 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2462 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2461 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2460 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2459 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2458 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2457 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2456 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2455 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2454 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2453 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2452 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2451 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2450 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2449 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2448 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2447 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2446 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2445 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2444 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2443 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2442 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2441 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2440 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2439 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2438 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2437 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2436 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2435 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2434 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2433 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2432 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2431 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2430 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2429 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2428 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2427 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2426 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2425 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2424 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2423 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2422 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2421 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2420 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2419 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2418 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2417 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2416 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2415 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2414 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2413 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2412 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2411 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2410 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2409 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2408 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2407 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2406 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2405 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2404 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2403 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2402 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2401 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_18 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_74 UIV ( .A(n1), .Y(SB) );
  ND2_2400 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2399 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2398 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2397 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2396 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2395 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2394 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2393 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2392 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2391 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2390 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2389 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2388 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2387 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2386 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2385 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2384 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2383 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2382 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2381 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2380 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2379 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2378 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2377 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2376 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2375 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2374 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2373 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2372 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2371 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2370 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2369 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2368 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2367 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2366 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2365 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2364 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2363 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2362 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2361 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2360 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2359 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2358 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2357 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2356 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2355 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2354 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2353 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2352 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2351 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2350 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2349 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2348 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2347 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2346 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2345 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2344 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2343 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2342 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2341 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2340 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2339 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2338 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2337 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2336 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2335 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2334 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2333 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2332 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2331 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2330 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2329 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2328 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2327 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2326 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2325 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2324 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2323 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2322 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2321 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2320 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2319 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2318 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2317 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2316 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2315 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2314 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2313 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2312 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2311 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2310 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2309 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2308 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2307 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2306 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2305 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_17 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_73 UIV ( .A(n1), .Y(SB) );
  ND2_2304 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2303 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2302 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2301 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2300 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2299 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2298 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2297 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2296 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2295 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2294 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2293 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2292 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2291 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2290 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2289 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2288 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2287 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2286 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2285 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2284 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2283 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2282 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2281 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2280 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2279 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2278 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2277 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2276 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2275 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2274 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2273 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2272 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2271 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2270 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2269 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2268 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2267 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2266 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2265 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2264 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2263 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2262 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2261 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2260 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2259 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2258 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2257 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2256 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2255 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2254 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2253 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2252 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2251 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2250 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2249 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2248 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2247 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2246 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2245 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2244 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2243 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2242 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2241 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2240 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2239 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2238 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2237 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2236 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2235 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2234 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2233 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2232 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2231 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2230 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2229 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2228 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2227 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2226 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2225 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2224 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2223 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2222 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2221 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2220 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2219 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2218 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2217 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2216 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2215 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2214 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2213 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2212 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2211 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2210 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2209 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_16 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_72 UIV ( .A(n1), .Y(SB) );
  ND2_2208 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2207 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2206 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2205 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2204 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2203 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2202 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2201 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2200 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2199 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2198 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2197 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2196 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2195 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2194 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2193 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2192 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2191 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2190 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2189 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2188 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2187 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2186 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2185 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2184 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2183 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2182 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2181 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2180 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2179 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2178 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2177 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2176 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2175 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2174 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2173 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2172 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2171 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2170 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2169 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2168 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2167 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2166 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2165 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2164 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2163 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2162 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2161 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2160 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2159 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2158 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2157 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2156 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2155 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2154 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2153 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2152 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2151 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2150 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2149 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2148 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2147 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2146 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2145 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2144 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2143 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2142 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2141 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2140 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2139 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2138 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2137 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2136 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2135 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2134 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2133 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2132 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2131 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2130 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2129 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2128 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2127 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2126 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2125 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2124 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2123 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2122 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2121 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2120 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2119 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2118 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2117 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2116 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2115 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2114 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2113 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_15 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_71 UIV ( .A(n1), .Y(SB) );
  ND2_2112 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2111 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2110 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2109 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2108 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2107 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2106 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2105 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2104 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2103 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2102 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2101 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2100 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2099 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2098 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2097 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2096 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_2095 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_2094 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_2093 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_2092 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_2091 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_2090 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_2089 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_2088 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_2087 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_2086 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_2085 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_2084 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_2083 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_2082 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_2081 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_2080 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_2079 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_2078 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_2077 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_2076 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_2075 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_2074 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_2073 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_2072 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_2071 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_2070 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_2069 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_2068 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_2067 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_2066 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_2065 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_2064 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_2063 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_2062 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_2061 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_2060 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_2059 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_2058 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_2057 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_2056 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_2055 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_2054 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_2053 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_2052 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_2051 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_2050 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_2049 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_2048 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_2047 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_2046 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_2045 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_2044 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_2043 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_2042 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_2041 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_2040 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_2039 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_2038 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_2037 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_2036 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_2035 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_2034 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_2033 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_2032 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_2031 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_2030 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_2029 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_2028 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_2027 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_2026 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_2025 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_2024 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_2023 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_2022 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_2021 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_2020 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_2019 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2018 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_2017 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_14 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_70 UIV ( .A(n1), .Y(SB) );
  ND2_2016 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_2015 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_2014 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_2013 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_2012 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_2011 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_2010 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_2009 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_2008 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_2007 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_2006 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_2005 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_2004 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_2003 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_2002 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_2001 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_2000 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1999 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1998 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1997 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1996 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1995 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1994 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1993 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1992 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1991 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1990 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1989 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1988 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1987 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1986 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1985 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1984 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1983 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1982 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1981 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1980 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1979 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1978 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1977 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1976 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1975 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1974 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1973 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1972 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1971 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1970 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1969 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1968 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1967 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1966 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1965 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1964 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1963 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1962 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1961 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1960 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1959 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1958 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1957 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1956 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1955 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1954 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1953 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1952 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1951 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1950 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1949 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1948 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1947 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1946 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1945 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1944 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1943 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1942 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1941 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1940 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1939 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1938 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1937 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1936 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1935 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1934 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1933 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1932 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1931 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1930 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1929 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1928 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1927 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1926 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1925 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1924 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1923 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1922 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1921 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_13 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_69 UIV ( .A(n1), .Y(SB) );
  ND2_1920 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1919 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1918 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1917 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1916 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1915 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1914 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1913 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1912 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1911 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1910 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1909 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1908 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1907 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1906 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1905 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1904 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1903 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1902 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1901 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1900 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1899 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1898 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1897 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1896 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1895 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1894 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1893 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1892 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1891 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1890 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1889 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1888 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1887 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1886 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1885 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1884 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1883 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1882 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1881 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1880 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1879 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1878 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1877 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1876 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1875 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1874 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1873 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1872 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1871 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1870 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1869 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1868 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1867 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1866 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1865 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1864 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1863 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1862 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1861 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1860 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1859 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1858 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1857 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1856 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1855 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1854 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1853 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1852 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1851 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1850 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1849 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1848 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1847 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1846 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1845 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1844 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1843 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1842 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1841 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1840 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1839 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1838 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1837 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1836 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1835 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1834 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1833 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1832 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1831 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1830 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1829 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1828 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1827 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1826 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1825 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_12 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_68 UIV ( .A(n1), .Y(SB) );
  ND2_1824 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1823 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1822 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1821 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1820 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1819 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1818 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1817 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1816 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1815 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1814 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1813 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1812 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1811 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1810 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1809 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1808 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1807 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1806 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1805 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1804 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1803 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1802 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1801 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1800 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1799 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1798 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1797 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1796 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1795 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1794 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1793 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1792 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1791 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1790 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1789 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1788 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1787 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1786 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1785 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1784 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1783 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1782 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1781 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1780 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1779 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1778 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1777 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1776 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1775 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1774 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1773 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1772 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1771 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1770 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1769 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1768 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1767 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1766 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1765 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1764 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1763 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1762 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1761 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1760 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1759 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1758 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1757 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1756 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1755 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1754 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1753 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1752 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1751 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1750 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1749 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1748 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1747 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1746 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1745 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1744 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1743 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1742 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1741 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1740 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1739 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1738 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1737 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1736 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1735 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1734 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1733 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1732 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1731 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1730 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1729 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_11 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_67 UIV ( .A(n1), .Y(SB) );
  ND2_1728 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1727 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1726 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1725 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1724 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1723 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1722 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1721 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1720 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1719 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1718 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1717 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1716 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1715 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1714 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1713 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1712 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1711 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1710 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1709 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1708 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1707 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1706 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1705 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1704 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1703 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1702 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1701 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1700 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1699 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1698 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1697 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1696 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1695 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1694 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1693 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1692 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1691 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1690 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1689 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1688 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1687 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1686 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1685 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1684 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1683 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1682 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1681 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1680 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1679 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1678 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1677 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1676 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1675 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1674 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1673 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1672 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1671 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1670 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1669 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1668 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1667 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1666 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1665 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1664 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1663 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1662 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1661 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1660 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1659 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1658 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1657 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1656 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1655 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1654 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1653 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1652 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1651 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1650 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1649 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1648 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1647 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1646 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1645 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1644 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1643 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1642 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1641 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1640 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1639 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1638 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1637 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1636 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1635 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1634 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1633 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_10 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_66 UIV ( .A(n1), .Y(SB) );
  ND2_1632 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1631 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1630 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1629 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1628 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1627 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1626 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1625 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1624 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1623 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1622 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1621 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1620 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1619 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1618 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1617 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1616 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1615 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1614 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1613 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1612 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1611 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1610 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1609 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1608 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1607 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1606 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1605 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1604 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1603 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1602 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1601 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1600 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1599 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1598 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1597 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1596 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1595 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1594 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1593 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1592 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1591 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1590 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1589 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1588 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1587 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1586 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1585 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1584 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1583 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1582 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1581 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1580 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1579 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1578 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1577 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1576 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1575 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1574 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1573 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1572 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1571 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1570 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1569 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1568 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1567 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1566 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1565 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1564 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1563 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1562 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1561 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1560 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1559 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1558 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1557 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1556 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1555 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1554 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1553 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1552 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1551 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1550 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1549 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1548 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1547 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1546 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1545 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1544 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1543 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1542 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1541 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1540 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1539 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1538 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1537 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_9 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_65 UIV ( .A(n1), .Y(SB) );
  ND2_1536 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1535 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1534 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1533 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1532 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1531 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1530 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1529 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1528 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1527 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1526 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1525 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1524 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1523 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1522 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1521 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1520 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1519 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1518 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1517 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1516 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1515 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1514 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1513 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1512 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1511 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1510 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1509 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1508 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1507 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1506 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1505 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1504 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1503 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1502 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1501 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1500 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1499 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1498 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1497 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1496 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1495 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1494 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1493 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1492 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1491 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1490 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1489 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1488 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1487 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1486 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1485 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1484 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1483 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1482 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1481 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1480 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1479 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1478 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1477 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1476 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1475 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1474 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1473 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1472 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1471 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1470 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1469 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1468 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1467 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1466 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1465 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1464 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1463 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1462 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1461 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1460 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1459 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1458 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1457 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1456 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1455 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1454 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1453 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1452 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1451 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1450 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1449 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1448 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1447 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1446 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1445 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1444 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1443 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1442 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1441 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_8 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_64 UIV ( .A(n1), .Y(SB) );
  ND2_1440 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1439 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1438 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1437 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1436 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1435 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1434 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1433 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1432 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1431 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1430 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1429 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1428 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1427 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1426 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1425 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1424 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1423 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1422 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1421 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1420 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1419 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1418 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1417 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1416 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1415 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1414 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1413 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1412 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1411 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1410 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1409 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1408 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1407 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1406 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1405 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1404 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1403 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1402 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1401 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1400 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1399 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1398 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1397 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1396 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1395 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1394 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1393 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1392 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1391 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1390 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1389 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1388 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1387 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1386 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1385 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1384 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1383 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1382 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1381 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1380 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1379 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1378 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1377 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1376 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1375 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1374 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1373 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1372 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1371 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1370 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1369 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1368 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1367 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1366 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1365 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1364 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1363 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1362 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1361 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1360 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1359 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1358 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1357 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1356 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1355 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1354 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1353 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1352 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1351 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1350 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1349 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1348 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1347 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1346 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1345 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_7 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_63 UIV ( .A(n1), .Y(SB) );
  ND2_1344 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1343 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1342 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1341 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1340 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1339 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1338 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1337 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1336 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1335 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1334 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1333 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1332 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1331 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1330 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1329 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1328 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1327 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1326 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1325 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1324 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1323 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1322 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1321 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1320 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1319 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1318 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1317 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1316 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1315 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1314 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1313 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1312 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1311 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1310 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1309 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1308 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1307 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1306 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1305 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1304 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1303 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1302 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1301 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1300 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1299 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1298 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1297 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1296 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1295 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1294 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1293 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1292 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1291 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1290 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1289 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1288 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1287 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1286 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1285 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1284 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1283 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1282 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1281 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1280 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1279 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1278 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1277 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1276 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1275 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1274 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1273 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1272 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1271 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1270 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1269 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1268 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1267 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1266 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1265 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1264 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1263 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1262 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1261 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1260 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1259 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1258 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1257 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1256 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1255 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1254 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1253 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1252 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1251 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1250 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1249 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_62 UIV ( .A(n1), .Y(SB) );
  ND2_1248 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1247 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1246 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1245 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1244 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1243 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1242 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1241 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1240 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1239 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1238 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1237 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1236 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1235 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1234 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1233 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1232 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1231 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1230 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1229 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1228 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1227 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1226 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1225 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1224 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1223 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1222 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1221 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1220 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1219 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1218 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1217 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1216 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1215 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1214 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1213 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1212 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1211 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1210 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1209 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1208 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1207 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1206 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1205 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1204 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1203 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1202 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1201 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1200 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1199 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1198 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1197 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1196 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1195 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1194 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1193 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1192 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1191 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1190 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1189 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1188 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1187 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1186 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1185 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1184 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1183 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1182 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1181 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1180 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1179 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1178 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1177 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1176 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1175 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1174 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1173 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1172 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1171 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1170 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1169 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1168 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1167 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1166 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1165 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1164 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1163 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1162 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1161 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1160 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1159 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1158 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1157 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1156 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1155 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1154 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1153 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_61 UIV ( .A(n1), .Y(SB) );
  ND2_1152 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1151 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1150 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1149 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1148 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1147 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1146 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1145 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1144 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1143 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1142 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1141 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1140 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1139 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1138 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1137 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1136 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1135 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1134 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1133 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1132 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1131 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1130 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1129 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1128 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1127 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1126 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1125 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1124 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1123 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1122 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1121 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1120 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1119 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1118 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1117 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1116 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1115 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1114 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1113 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1112 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1111 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1110 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1109 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1108 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1107 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1106 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1105 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1104 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1103 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1102 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1101 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1100 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1099 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1098 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1097 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1096 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_1095 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_1094 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_1093 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_1092 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_1091 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_1090 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_1089 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_1088 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_1087 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_1086 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_1085 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_1084 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_1083 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_1082 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_1081 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_1080 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_1079 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_1078 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_1077 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_1076 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_1075 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_1074 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_1073 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_1072 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_1071 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_1070 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_1069 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_1068 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_1067 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_1066 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_1065 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_1064 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_1063 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_1062 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_1061 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_1060 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_1059 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_1058 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_1057 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_60 UIV ( .A(n1), .Y(SB) );
  ND2_1056 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_1055 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_1054 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_1053 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_1052 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_1051 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_1050 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_1049 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_1048 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_1047 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_1046 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_1045 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_1044 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_1043 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_1042 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_1041 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_1040 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_1039 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_1038 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_1037 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_1036 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_1035 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_1034 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_1033 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_1032 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_1031 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_1030 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_1029 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_1028 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_1027 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_1026 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_1025 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_1024 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_1023 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_1022 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_1021 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_1020 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_1019 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_1018 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_1017 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_1016 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_1015 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_1014 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_1013 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_1012 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_1011 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_1010 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_1009 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_1008 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_1007 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_1006 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_1005 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_1004 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_1003 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_1002 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_1001 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_1000 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_999 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_998 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_997 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_996 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_995 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_994 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_993 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_992 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_991 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_990 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_989 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_988 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_987 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_986 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_985 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_984 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_983 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_982 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_981 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_980 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_979 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_978 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_977 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_976 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_975 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_974 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_973 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_972 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_971 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_970 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_969 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_968 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_967 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_966 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_965 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_964 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_963 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_962 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_961 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_59 UIV ( .A(n1), .Y(SB) );
  ND2_960 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_959 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_958 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_957 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_956 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_955 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_954 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_953 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_952 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_951 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_950 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_949 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_948 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_947 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_946 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_945 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_944 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_943 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_942 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_941 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_940 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_939 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_938 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_937 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_936 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_935 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_934 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_933 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_932 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_931 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_930 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_929 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_928 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_927 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_926 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_925 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_924 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_923 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_922 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_921 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_920 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_919 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_918 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_917 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_916 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_915 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_914 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_913 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_912 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_911 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_910 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_909 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_908 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_907 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_906 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_905 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_904 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_903 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_902 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_901 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_900 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_899 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_898 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_897 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_896 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_895 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_894 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_893 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_892 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_891 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_890 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_889 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_888 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_887 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_886 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_885 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_884 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_883 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_882 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_881 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_880 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_879 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_878 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_877 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_876 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_875 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_874 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_873 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_872 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_871 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_870 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_869 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_868 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_867 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_866 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_865 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_58 UIV ( .A(n1), .Y(SB) );
  ND2_864 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_863 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_862 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_861 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_860 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_859 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_858 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_857 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_856 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_855 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_854 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_853 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_852 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_851 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_850 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_849 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_848 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_847 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_846 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_845 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_844 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_843 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_842 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_841 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_840 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_839 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_838 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_837 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_836 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_835 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_834 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_833 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_832 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_831 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_830 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_829 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_828 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_827 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_826 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_825 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_824 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_823 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_822 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_821 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_820 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_819 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_818 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_817 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_816 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_815 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_814 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_813 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_812 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_811 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_810 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_809 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_808 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_807 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_806 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_805 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_804 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_803 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_802 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_801 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_800 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_799 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_798 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_797 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_796 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_795 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_794 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_793 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_792 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_791 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_790 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_789 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_788 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_787 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_786 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_785 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_784 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_783 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_782 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_781 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_780 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_779 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_778 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_777 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_776 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_775 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_774 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_773 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_772 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_771 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_770 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_769 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GENERIC_N32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_57 UIV ( .A(n1), .Y(SB) );
  ND2_768 UND1_31 ( .A(A[31]), .B(n3), .Y(Y1[31]) );
  ND2_767 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_766 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_765 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_764 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_763 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_762 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_761 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_760 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_759 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_758 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_757 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_756 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_755 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_754 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_753 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_752 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_751 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_750 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_749 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_748 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_747 UND1_24 ( .A(A[24]), .B(n2), .Y(Y1[24]) );
  ND2_746 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_745 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_744 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_743 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_742 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_741 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_740 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_739 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_738 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_737 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_736 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_735 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_734 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_733 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_732 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_731 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_730 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_729 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_728 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_727 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_726 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_725 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_724 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_723 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_722 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_721 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_720 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_719 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_718 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_717 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_716 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_715 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_714 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_713 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_712 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_711 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_710 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_709 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_708 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  ND2_707 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_706 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_705 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_704 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_703 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_702 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_701 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_700 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_699 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_698 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_697 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_696 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_695 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_694 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_693 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_692 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_691 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_690 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_689 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_688 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_687 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_686 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_685 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_684 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_683 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_682 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_681 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_680 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_679 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_678 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_677 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_676 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_675 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_674 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_673 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module P4adder_N32_PowerN5_6 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;

  wire   [7:0] sCout;

  sparce_tree_POWER5_6 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_6 USum_generator ( .A(A), .B(B), .Ci(sCout), 
        .S(S) );
endmodule


module P4adder_N32_PowerN5_5 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;
  wire   n1, n2;
  wire   [7:0] sCout;

  sparce_tree_POWER5_5 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_5 USum_generator ( .A(A), .B({B[31:20], n2, 
        B[18:0]}), .Ci(sCout), .S(S) );
  INV_X1 U1 ( .A(B[19]), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
endmodule


module P4adder_N32_PowerN5_4 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;

  wire   [7:0] sCout;

  sparce_tree_POWER5_4 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_4 USum_generator ( .A(A), .B(B), .Ci(sCout), 
        .S(S) );
endmodule


module P4adder_N32_PowerN5_3 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;

  wire   [7:0] sCout;

  sparce_tree_POWER5_3 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_3 USum_generator ( .A(A), .B(B), .Ci(sCout), 
        .S(S) );
endmodule


module P4adder_N32_PowerN5_2 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;
  wire   n1, n2, n3;
  wire   [7:0] sCout;

  sparce_tree_POWER5_2 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_2 USum_generator ( .A(A), .B({B[31:28], n3, 
        B[26:24], n2, B[22:0]}), .Ci(sCout), .S(S) );
  INV_X1 U1 ( .A(B[23]), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
  CLKBUF_X1 U3 ( .A(B[27]), .Z(n3) );
endmodule


module P4adder_N32_PowerN5_1 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;

  wire   [7:0] sCout;

  sparce_tree_POWER5_1 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_1 USum_generator ( .A(A), .B(B), .Ci(sCout), 
        .S(S) );
endmodule


module booth_mux_generic_N32_7 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  MUX21_GENERIC_N32_28 mux1 ( .A(A_neg), .B(A), .SEL(n3), .Y(mux_A) );
  MUX21_GENERIC_N32_27 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n3), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_26 mux3 ( .A(mux_2a), .B(Zero), .SEL(n1), .Y(mux_zero_2a)
         );
  MUX21_GENERIC_N32_25 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(n2), .Y(Y) );
  BUF_X1 U1 ( .A(SEL[2]), .Z(n3) );
  XOR2_X1 U2 ( .A(n3), .B(SEL[1]), .Z(n1) );
  XOR2_X1 U3 ( .A(SEL[1]), .B(SEL[0]), .Z(n2) );
endmodule


module booth_mux_generic_N32_6 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   selmux3, n1, n2;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  XOR2_X1 U2 ( .A(n2), .B(SEL[1]), .Z(selmux3) );
  MUX21_GENERIC_N32_24 mux1 ( .A(A_neg), .B(A), .SEL(n2), .Y(mux_A) );
  MUX21_GENERIC_N32_23 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n2), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_22 mux3 ( .A(mux_2a), .B(Zero), .SEL(selmux3), .Y(
        mux_zero_2a) );
  MUX21_GENERIC_N32_21 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(n1), .Y(Y) );
  XOR2_X1 U1 ( .A(SEL[1]), .B(SEL[0]), .Z(n1) );
  BUF_X1 U3 ( .A(SEL[2]), .Z(n2) );
endmodule


module booth_mux_generic_N32_5 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   selmux3, selmux4, n1;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  XOR2_X1 U1 ( .A(SEL[1]), .B(SEL[0]), .Z(selmux4) );
  XOR2_X1 U2 ( .A(n1), .B(SEL[1]), .Z(selmux3) );
  MUX21_GENERIC_N32_20 mux1 ( .A(A_neg), .B(A), .SEL(n1), .Y(mux_A) );
  MUX21_GENERIC_N32_19 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n1), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_18 mux3 ( .A(mux_2a), .B(Zero), .SEL(selmux3), .Y(
        mux_zero_2a) );
  MUX21_GENERIC_N32_17 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(selmux4), .Y(Y)
         );
  BUF_X1 U3 ( .A(SEL[2]), .Z(n1) );
endmodule


module booth_mux_generic_N32_4 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   selmux3, selmux4, n1;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  XOR2_X1 U1 ( .A(SEL[1]), .B(SEL[0]), .Z(selmux4) );
  XOR2_X1 U2 ( .A(n1), .B(SEL[1]), .Z(selmux3) );
  MUX21_GENERIC_N32_16 mux1 ( .A(A_neg), .B(A), .SEL(n1), .Y(mux_A) );
  MUX21_GENERIC_N32_15 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n1), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_14 mux3 ( .A(mux_2a), .B(Zero), .SEL(selmux3), .Y(
        mux_zero_2a) );
  MUX21_GENERIC_N32_13 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(selmux4), .Y(Y)
         );
  BUF_X1 U3 ( .A(SEL[2]), .Z(n1) );
endmodule


module booth_mux_generic_N32_3 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   selmux3, selmux4, n1;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  XOR2_X1 U1 ( .A(SEL[1]), .B(SEL[0]), .Z(selmux4) );
  XOR2_X1 U2 ( .A(n1), .B(SEL[1]), .Z(selmux3) );
  MUX21_GENERIC_N32_12 mux1 ( .A(A_neg), .B(A), .SEL(n1), .Y(mux_A) );
  MUX21_GENERIC_N32_11 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n1), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_10 mux3 ( .A(mux_2a), .B(Zero), .SEL(selmux3), .Y(
        mux_zero_2a) );
  MUX21_GENERIC_N32_9 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(selmux4), .Y(Y)
         );
  BUF_X1 U3 ( .A(SEL[2]), .Z(n1) );
endmodule


module booth_mux_generic_N32_2 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   selmux3, selmux4, n1;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  XOR2_X1 U1 ( .A(SEL[1]), .B(SEL[0]), .Z(selmux4) );
  XOR2_X1 U2 ( .A(n1), .B(SEL[1]), .Z(selmux3) );
  MUX21_GENERIC_N32_8 mux1 ( .A(A_neg), .B(A), .SEL(n1), .Y(mux_A) );
  MUX21_GENERIC_N32_7 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n1), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_6 mux3 ( .A(mux_2a), .B(Zero), .SEL(selmux3), .Y(
        mux_zero_2a) );
  MUX21_GENERIC_N32_5 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(selmux4), .Y(Y)
         );
  BUF_X1 U3 ( .A(SEL[2]), .Z(n1) );
endmodule


module booth_mux_generic_N32_1 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   selmux3, selmux4, n1;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  XOR2_X1 U1 ( .A(SEL[1]), .B(SEL[0]), .Z(selmux4) );
  XOR2_X1 U2 ( .A(n1), .B(SEL[1]), .Z(selmux3) );
  MUX21_GENERIC_N32_4 mux1 ( .A(A_neg), .B(A), .SEL(n1), .Y(mux_A) );
  MUX21_GENERIC_N32_3 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n1), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_2 mux3 ( .A(mux_2a), .B(Zero), .SEL(selmux3), .Y(
        mux_zero_2a) );
  MUX21_GENERIC_N32_1 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(selmux4), .Y(Y)
         );
  BUF_X1 U3 ( .A(SEL[2]), .Z(n1) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_GENERIC_N4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_56 UIV ( .A(SEL), .Y(SB) );
  ND2_672 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_671 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_670 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_669 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_668 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_667 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_666 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_665 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_664 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_663 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_662 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_661 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module RCA_generic_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_447 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_446 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_445 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module cs_generic_N4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_0 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_111 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_0 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module block_pg_0 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n2;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n2) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n2), .ZN(Gij) );
endmodule


module block_g_0 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n2) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module Sum_generator_Nbit32_Nblock8_0 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_0 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  cs_generic_N4_55 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4])
         );
  cs_generic_N4_54 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  cs_generic_N4_53 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_52 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_51 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_50 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_49 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sparce_tree_POWER5_0 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, p1, g1, \matrixG[16][16] , \matrixG[16][15] , \matrixG[16][13] ,
         \matrixG[16][9] , \matrixG[15][15] , \matrixG[14][14] ,
         \matrixG[14][13] , \matrixG[13][13] , \matrixG[12][12] ,
         \matrixG[12][11] , \matrixG[12][9] , \matrixG[11][11] ,
         \matrixG[10][10] , \matrixG[10][9] , \matrixG[9][9] , \matrixG[8][8] ,
         \matrixG[8][7] , \matrixG[8][5] , \matrixG[7][7] , \matrixG[6][6] ,
         \matrixG[6][5] , \matrixG[5][5] , \matrixG[4][4] , \matrixG[4][3] ,
         \matrixG[3][3] , \matrixG[2][2] , \matrixG[2][1] , \matrixG[1][1] ,
         \matrixP[16][16] , \matrixP[16][15] , \matrixP[16][13] ,
         \matrixP[16][9] , \matrixP[15][15] , \matrixP[14][14] ,
         \matrixP[14][13] , \matrixP[13][13] , \matrixP[12][12] ,
         \matrixP[12][11] , \matrixP[12][9] , \matrixP[11][11] ,
         \matrixP[10][10] , \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] ,
         \matrixP[8][7] , \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] ,
         \matrixP[6][5] , \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] ,
         \matrixP[3][3] , \matrixP[2][2] , \matrixP[32][32] ,
         \matrixP[32][31] , \matrixP[32][29] , \matrixP[32][25] ,
         \matrixP[32][17] , \matrixP[31][31] , \matrixP[30][30] ,
         \matrixP[30][29] , \matrixP[29][29] , \matrixP[28][28] ,
         \matrixP[28][27] , \matrixP[28][25] , \matrixP[28][17] ,
         \matrixP[27][27] , \matrixP[26][26] , \matrixP[26][25] ,
         \matrixP[25][25] , \matrixP[24][24] , \matrixP[24][23] ,
         \matrixP[24][21] , \matrixP[24][17] , \matrixP[23][23] ,
         \matrixP[22][22] , \matrixP[22][21] , \matrixP[21][21] ,
         \matrixP[20][20] , \matrixP[20][19] , \matrixP[20][17] ,
         \matrixP[19][19] , \matrixP[18][18] , \matrixP[18][17] ,
         \matrixP[17][17] , \matrixG[32][32] , \matrixG[32][31] ,
         \matrixG[32][29] , \matrixG[32][25] , \matrixG[32][17] ,
         \matrixG[31][31] , \matrixG[30][30] , \matrixG[30][29] ,
         \matrixG[29][29] , \matrixG[28][28] , \matrixG[28][27] ,
         \matrixG[28][25] , \matrixG[28][17] , \matrixG[27][27] ,
         \matrixG[26][26] , \matrixG[26][25] , \matrixG[25][25] ,
         \matrixG[24][24] , \matrixG[24][23] , \matrixG[24][21] ,
         \matrixG[24][17] , \matrixG[23][23] , \matrixG[22][22] ,
         \matrixG[22][21] , \matrixG[21][21] , \matrixG[20][20] ,
         \matrixG[20][19] , \matrixG[20][17] , \matrixG[19][19] ,
         \matrixG[18][18] , \matrixG[18][17] , \matrixG[17][17] ;
  assign Cout[0] = Ci;

  XOR2_X1 U33 ( .A(B[1]), .B(A[1]), .Z(p1) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U46 ( .A(B[28]), .B(A[28]), .Z(\matrixP[28][28] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U50 ( .A(B[24]), .B(A[24]), .Z(\matrixP[24][24] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U54 ( .A(B[20]), .B(A[20]), .Z(\matrixP[20][20] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  block_g_0 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_69 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_0 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), .Gik(
        \matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), .Gij(
        \matrixG[4][3] ) );
  block_pg_188 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), 
        .Gik(\matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), 
        .Gij(\matrixG[6][5] ) );
  block_pg_187 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), 
        .Gik(\matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), 
        .Gij(\matrixG[8][7] ) );
  block_pg_186 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_185 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_184 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_183 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_182 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_181 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_180 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_179 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_178 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_177 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_176 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_175 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_68 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(Cout[1]) );
  block_pg_174 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), 
        .Gik(\matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), 
        .Gij(\matrixG[8][5] ) );
  block_pg_173 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_172 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_171 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_170 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_169 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_168 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_67 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(
        Cout[1]), .Gij(Cout[2]) );
  block_pg_167 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_166 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_165 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_66 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[4]) );
  block_g_65 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(Cout[2]), .Gij(Cout[3]) );
  block_pg_164 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_163 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_64 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_63 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[7]) );
  block_g_62 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[6]) );
  block_g_61 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[5]) );
  XOR2_X2 U1 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  AND2_X1 U2 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  XOR2_X1 U3 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  AND2_X1 U4 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U5 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U6 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U7 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U8 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U9 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  AND2_X1 U10 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U11 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  AND2_X1 U12 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
  AND2_X1 U13 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U14 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  AND2_X1 U15 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  AND2_X1 U16 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U17 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U18 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U19 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U20 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U21 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U22 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U23 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U24 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  AND2_X1 U25 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U26 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U27 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U28 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U29 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U30 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U31 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  AND2_X1 U32 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U58 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U62 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
endmodule


module MUX21_GENERIC_N32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  IV_0 UIV ( .A(n1), .Y(SB) );
  ND2_0 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  ND2_3743 UND2_31 ( .A(B[31]), .B(n6), .Y(Y2[31]) );
  ND2_3742 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  ND2_3741 UND1_30 ( .A(A[30]), .B(n3), .Y(Y1[30]) );
  ND2_3740 UND2_30 ( .A(B[30]), .B(n6), .Y(Y2[30]) );
  ND2_3739 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  ND2_3738 UND1_29 ( .A(A[29]), .B(n3), .Y(Y1[29]) );
  ND2_3737 UND2_29 ( .A(B[29]), .B(n6), .Y(Y2[29]) );
  ND2_3736 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  ND2_3735 UND1_28 ( .A(A[28]), .B(n3), .Y(Y1[28]) );
  ND2_3734 UND2_28 ( .A(B[28]), .B(n6), .Y(Y2[28]) );
  ND2_3733 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  ND2_3732 UND1_27 ( .A(A[27]), .B(n3), .Y(Y1[27]) );
  ND2_3731 UND2_27 ( .A(B[27]), .B(n6), .Y(Y2[27]) );
  ND2_3730 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  ND2_3729 UND1_26 ( .A(A[26]), .B(n3), .Y(Y1[26]) );
  ND2_3728 UND2_26 ( .A(B[26]), .B(n6), .Y(Y2[26]) );
  ND2_3727 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  ND2_3726 UND1_25 ( .A(A[25]), .B(n3), .Y(Y1[25]) );
  ND2_3725 UND2_25 ( .A(B[25]), .B(n5), .Y(Y2[25]) );
  ND2_3724 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  ND2_3723 UND1_24 ( .A(A[24]), .B(n3), .Y(Y1[24]) );
  ND2_3722 UND2_24 ( .A(B[24]), .B(n5), .Y(Y2[24]) );
  ND2_3721 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  ND2_3720 UND1_23 ( .A(A[23]), .B(n2), .Y(Y1[23]) );
  ND2_3719 UND2_23 ( .A(B[23]), .B(n5), .Y(Y2[23]) );
  ND2_3718 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  ND2_3717 UND1_22 ( .A(A[22]), .B(n2), .Y(Y1[22]) );
  ND2_3716 UND2_22 ( .A(B[22]), .B(n5), .Y(Y2[22]) );
  ND2_3715 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  ND2_3714 UND1_21 ( .A(A[21]), .B(n2), .Y(Y1[21]) );
  ND2_3713 UND2_21 ( .A(B[21]), .B(n5), .Y(Y2[21]) );
  ND2_3712 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  ND2_3711 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  ND2_3710 UND2_20 ( .A(B[20]), .B(n5), .Y(Y2[20]) );
  ND2_3709 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  ND2_3708 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  ND2_3707 UND2_19 ( .A(B[19]), .B(n5), .Y(Y2[19]) );
  ND2_3706 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  ND2_3705 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  ND2_3704 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  ND2_3703 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  ND2_3702 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  ND2_3701 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  ND2_3700 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  ND2_3699 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  ND2_3698 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  ND2_3697 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  ND2_3696 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  ND2_3695 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  ND2_3694 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  ND2_3693 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  ND2_3692 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  ND2_3691 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  ND2_3690 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  ND2_3689 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  ND2_3688 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  ND2_3687 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  ND2_3686 UND2_12 ( .A(B[12]), .B(n4), .Y(Y2[12]) );
  ND2_3685 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  ND2_3684 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  ND2_3683 UND2_11 ( .A(B[11]), .B(n4), .Y(Y2[11]) );
  ND2_3682 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  ND2_3681 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  ND2_3680 UND2_10 ( .A(B[10]), .B(n4), .Y(Y2[10]) );
  ND2_3679 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  ND2_3678 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  ND2_3677 UND2_9 ( .A(B[9]), .B(n4), .Y(Y2[9]) );
  ND2_3676 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  ND2_3675 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  ND2_3674 UND2_8 ( .A(B[8]), .B(n4), .Y(Y2[8]) );
  ND2_3673 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  ND2_3672 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  ND2_3671 UND2_7 ( .A(B[7]), .B(n4), .Y(Y2[7]) );
  ND2_3670 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  ND2_3669 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  ND2_3668 UND2_6 ( .A(B[6]), .B(n4), .Y(Y2[6]) );
  ND2_3667 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  ND2_3666 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  ND2_3665 UND2_5 ( .A(B[5]), .B(n4), .Y(Y2[5]) );
  ND2_3664 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  ND2_3663 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  ND2_3662 UND2_4 ( .A(B[4]), .B(n4), .Y(Y2[4]) );
  ND2_3661 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  ND2_3660 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_3659 UND2_3 ( .A(B[3]), .B(n4), .Y(Y2[3]) );
  ND2_3658 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_3657 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_3656 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  ND2_3655 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_3654 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_3653 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  ND2_3652 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3651 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_3650 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  ND2_3649 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  CLKBUF_X1 U1 ( .A(SEL), .Z(n3) );
  CLKBUF_X1 U2 ( .A(SB), .Z(n6) );
  BUF_X1 U3 ( .A(SB), .Z(n4) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SB), .Z(n5) );
  BUF_X1 U6 ( .A(SEL), .Z(n2) );
endmodule


module P4adder_N32_PowerN5_0 ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;

  wire   [7:0] sCout;

  sparce_tree_POWER5_0 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, 
        sCout}) );
  Sum_generator_Nbit32_Nblock8_0 USum_generator ( .A(A), .B(B), .Ci(sCout), 
        .S(S) );
endmodule


module booth_mux_generic_N32_0 ( Zero, A, A_neg, A_double, A_neg_double, SEL, 
        Y );
  input [31:0] Zero;
  input [31:0] A;
  input [31:0] A_neg;
  input [31:0] A_double;
  input [31:0] A_neg_double;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3;
  wire   [31:0] mux_A;
  wire   [31:0] mux_2a;
  wire   [31:0] mux_zero_2a;

  MUX21_GENERIC_N32_0 mux1 ( .A(A_neg), .B(A), .SEL(n3), .Y(mux_A) );
  MUX21_GENERIC_N32_31 mux2 ( .A(A_neg_double), .B(A_double), .SEL(n3), .Y(
        mux_2a) );
  MUX21_GENERIC_N32_30 mux3 ( .A(mux_2a), .B(Zero), .SEL(n2), .Y(mux_zero_2a)
         );
  MUX21_GENERIC_N32_29 mux4 ( .A(mux_A), .B(mux_zero_2a), .SEL(n1), .Y(Y) );
  XOR2_X1 U1 ( .A(n3), .B(SEL[1]), .Z(n2) );
  XOR2_X1 U2 ( .A(SEL[1]), .B(SEL[0]), .Z(n1) );
  BUF_X4 U3 ( .A(SEL[2]), .Z(n3) );
endmodule


module boothmul_Nbit16 ( A, B, Res );
  input [15:0] A;
  input [15:0] B;
  output [31:0] Res;
  wire   N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13,
         \tmp_A_neg[7][31] , \tmp_A_neg[7][30] , \tmp_A_neg[7][29] ,
         \tmp_A_neg[7][28] , \tmp_A_neg[7][27] , \tmp_A_neg[7][26] ,
         \tmp_A_neg[7][25] , \tmp_A_neg[7][24] , \tmp_A_neg[7][23] ,
         \tmp_A_neg[7][22] , \tmp_A_neg[7][21] , \tmp_A_neg[7][20] ,
         \tmp_A_neg[7][19] , \tmp_A_neg[7][18] , \tmp_A_neg[7][17] ,
         \tmp_A_neg[7][16] , \tmp_A_neg[7][15] , \tmp_A_neg[6][31] ,
         \tmp_A_neg[6][30] , \tmp_A_neg[6][29] , \tmp_A_neg[6][28] ,
         \tmp_A_neg[6][27] , \tmp_A_neg[6][26] , \tmp_A_neg[6][25] ,
         \tmp_A_neg[6][24] , \tmp_A_neg[6][23] , \tmp_A_neg[6][22] ,
         \tmp_A_neg[6][21] , \tmp_A_neg[6][20] , \tmp_A_neg[6][19] ,
         \tmp_A_neg[6][18] , \tmp_A_neg[6][17] , \tmp_A_neg[6][16] ,
         \tmp_A_neg[6][15] , \tmp_A_neg[6][14] , \tmp_A_neg[6][13] ,
         \tmp_A_neg[5][31] , \tmp_A_neg[5][30] , \tmp_A_neg[5][29] ,
         \tmp_A_neg[5][28] , \tmp_A_neg[5][27] , \tmp_A_neg[5][26] ,
         \tmp_A_neg[5][25] , \tmp_A_neg[5][24] , \tmp_A_neg[5][23] ,
         \tmp_A_neg[5][22] , \tmp_A_neg[5][21] , \tmp_A_neg[5][20] ,
         \tmp_A_neg[5][19] , \tmp_A_neg[5][18] , \tmp_A_neg[5][17] ,
         \tmp_A_neg[5][16] , \tmp_A_neg[5][15] , \tmp_A_neg[5][14] ,
         \tmp_A_neg[5][13] , \tmp_A_neg[5][12] , \tmp_A_neg[5][11] ,
         \tmp_A_neg[5][10] , \tmp_A_neg[4][31] , \tmp_A_neg[4][23] ,
         \tmp_A_neg[4][22] , \tmp_A_neg[4][21] , \tmp_A_neg[4][20] ,
         \tmp_A_neg[4][19] , \tmp_A_neg[4][18] , \tmp_A_neg[4][17] ,
         \tmp_A_neg[4][16] , \tmp_A_neg[4][15] , \tmp_A_neg[4][14] ,
         \tmp_A_neg[4][13] , \tmp_A_neg[4][12] , \tmp_A_neg[4][11] ,
         \tmp_A_neg[4][10] , \tmp_A_neg[4][9] , \tmp_A_neg[3][31] ,
         \tmp_A_neg[3][21] , \tmp_A_neg[3][20] , \tmp_A_neg[3][19] ,
         \tmp_A_neg[3][18] , \tmp_A_neg[3][17] , \tmp_A_neg[3][16] ,
         \tmp_A_neg[3][15] , \tmp_A_neg[3][14] , \tmp_A_neg[3][13] ,
         \tmp_A_neg[3][12] , \tmp_A_neg[3][11] , \tmp_A_neg[3][10] ,
         \tmp_A_neg[3][9] , \tmp_A_neg[3][8] , \tmp_A_neg[3][7] ,
         \tmp_A_neg[2][31] , \tmp_A_neg[2][19] , \tmp_A_neg[2][18] ,
         \tmp_A_neg[2][17] , \tmp_A_neg[2][16] , \tmp_A_neg[2][15] ,
         \tmp_A_neg[2][14] , \tmp_A_neg[2][13] , \tmp_A_neg[2][12] ,
         \tmp_A_neg[2][11] , \tmp_A_neg[2][10] , \tmp_A_neg[2][9] ,
         \tmp_A_neg[2][8] , \tmp_A_neg[2][7] , \tmp_A_neg[2][6] ,
         \tmp_A_neg[2][5] , \tmp_A_neg[1][31] , \tmp_A_neg[1][17] ,
         \tmp_A_neg[1][16] , \tmp_A_neg[1][15] , \tmp_A_neg[1][14] ,
         \tmp_A_neg[1][13] , \tmp_A_neg[1][12] , \tmp_A_neg[1][11] ,
         \tmp_A_neg[1][10] , \tmp_A_neg[1][9] , \tmp_A_neg[1][8] ,
         \tmp_A_neg[1][7] , \tmp_A_neg[1][6] , \tmp_A_neg[1][5] ,
         \tmp_A_neg[1][4] , \tmp_A_neg[1][3] , \tmp_A_neg[0][31] ,
         \tmp_A_neg[0][15] , \tmp_A_neg[0][14] , \tmp_A_neg[0][13] ,
         \tmp_A_neg[0][12] , \tmp_A_neg[0][11] , \tmp_A_neg[0][10] ,
         \tmp_A_neg[0][9] , \tmp_A_neg[0][8] , \tmp_A_neg[0][7] ,
         \tmp_A_neg[0][6] , \tmp_A_neg[0][5] , \tmp_A_neg[0][4] ,
         \tmp_A_neg[0][3] , \tmp_A_neg[0][2] , \tmp_A_neg[0][1] ,
         \tmp_A_neg_double[7][31] , \tmp_A_neg_double[7][30] ,
         \tmp_A_neg_double[7][29] , \tmp_A_neg_double[7][28] ,
         \tmp_A_neg_double[7][27] , \tmp_A_neg_double[7][26] ,
         \tmp_A_neg_double[7][25] , \tmp_A_neg_double[7][24] ,
         \tmp_A_neg_double[7][23] , \tmp_A_neg_double[7][22] ,
         \tmp_A_neg_double[7][21] , \tmp_A_neg_double[7][20] ,
         \tmp_A_neg_double[7][19] , \tmp_A_neg_double[7][18] ,
         \tmp_A_neg_double[7][17] , \tmp_A_neg_double[7][16] ,
         \tmp_A_neg_double[6][31] , \tmp_A_neg_double[6][30] ,
         \tmp_A_neg_double[6][29] , \tmp_A_neg_double[6][28] ,
         \tmp_A_neg_double[6][27] , \tmp_A_neg_double[6][26] ,
         \tmp_A_neg_double[6][25] , \tmp_A_neg_double[6][24] ,
         \tmp_A_neg_double[6][23] , \tmp_A_neg_double[6][22] ,
         \tmp_A_neg_double[6][21] , \tmp_A_neg_double[6][20] ,
         \tmp_A_neg_double[6][19] , \tmp_A_neg_double[6][18] ,
         \tmp_A_neg_double[6][17] , \tmp_A_neg_double[6][16] ,
         \tmp_A_neg_double[6][15] , \tmp_A_neg_double[6][14] ,
         \tmp_A_neg_double[5][31] , \tmp_A_neg_double[5][30] ,
         \tmp_A_neg_double[5][29] , \tmp_A_neg_double[5][28] ,
         \tmp_A_neg_double[5][27] , \tmp_A_neg_double[5][26] ,
         \tmp_A_neg_double[5][25] , \tmp_A_neg_double[5][24] ,
         \tmp_A_neg_double[5][23] , \tmp_A_neg_double[5][22] ,
         \tmp_A_neg_double[5][21] , \tmp_A_neg_double[5][20] ,
         \tmp_A_neg_double[5][19] , \tmp_A_neg_double[5][18] ,
         \tmp_A_neg_double[5][17] , \tmp_A_neg_double[5][16] ,
         \tmp_A_neg_double[5][15] , \tmp_A_neg_double[5][14] ,
         \tmp_A_neg_double[5][13] , \tmp_A_neg_double[5][12] ,
         \tmp_A_neg_double[5][11] , \tmp_A_neg_double[4][31] ,
         \tmp_A_neg_double[4][24] , \tmp_A_neg_double[4][23] ,
         \tmp_A_neg_double[4][22] , \tmp_A_neg_double[4][21] ,
         \tmp_A_neg_double[4][20] , \tmp_A_neg_double[4][19] ,
         \tmp_A_neg_double[4][18] , \tmp_A_neg_double[4][17] ,
         \tmp_A_neg_double[4][16] , \tmp_A_neg_double[4][15] ,
         \tmp_A_neg_double[4][14] , \tmp_A_neg_double[4][13] ,
         \tmp_A_neg_double[4][12] , \tmp_A_neg_double[4][11] ,
         \tmp_A_neg_double[4][10] , \tmp_A_neg_double[3][31] ,
         \tmp_A_neg_double[3][22] , \tmp_A_neg_double[3][21] ,
         \tmp_A_neg_double[3][20] , \tmp_A_neg_double[3][19] ,
         \tmp_A_neg_double[3][18] , \tmp_A_neg_double[3][17] ,
         \tmp_A_neg_double[3][16] , \tmp_A_neg_double[3][15] ,
         \tmp_A_neg_double[3][14] , \tmp_A_neg_double[3][13] ,
         \tmp_A_neg_double[3][12] , \tmp_A_neg_double[3][11] ,
         \tmp_A_neg_double[3][10] , \tmp_A_neg_double[3][9] ,
         \tmp_A_neg_double[3][8] , \tmp_A_neg_double[2][31] ,
         \tmp_A_neg_double[2][20] , \tmp_A_neg_double[2][19] ,
         \tmp_A_neg_double[2][18] , \tmp_A_neg_double[2][17] ,
         \tmp_A_neg_double[2][16] , \tmp_A_neg_double[2][15] ,
         \tmp_A_neg_double[2][14] , \tmp_A_neg_double[2][13] ,
         \tmp_A_neg_double[2][12] , \tmp_A_neg_double[2][11] ,
         \tmp_A_neg_double[2][10] , \tmp_A_neg_double[2][9] ,
         \tmp_A_neg_double[2][8] , \tmp_A_neg_double[2][7] ,
         \tmp_A_neg_double[2][6] , \tmp_A_neg_double[1][31] ,
         \tmp_A_neg_double[1][18] , \tmp_A_neg_double[1][17] ,
         \tmp_A_neg_double[1][16] , \tmp_A_neg_double[1][15] ,
         \tmp_A_neg_double[1][14] , \tmp_A_neg_double[1][13] ,
         \tmp_A_neg_double[1][12] , \tmp_A_neg_double[1][11] ,
         \tmp_A_neg_double[1][10] , \tmp_A_neg_double[1][9] ,
         \tmp_A_neg_double[1][8] , \tmp_A_neg_double[1][7] ,
         \tmp_A_neg_double[1][6] , \tmp_A_neg_double[1][5] ,
         \tmp_A_neg_double[1][4] , \tmp_A_neg_double[0][31] ,
         \tmp_A_neg_double[0][16] , \tmp_A_neg_double[0][15] ,
         \tmp_A_neg_double[0][14] , \tmp_A_neg_double[0][13] ,
         \tmp_A_neg_double[0][12] , \tmp_A_neg_double[0][11] ,
         \tmp_A_neg_double[0][10] , \tmp_A_neg_double[0][9] ,
         \tmp_A_neg_double[0][8] , \tmp_A_neg_double[0][7] ,
         \tmp_A_neg_double[0][6] , \tmp_A_neg_double[0][5] ,
         \tmp_A_neg_double[0][4] , \tmp_A_neg_double[0][3] ,
         \tmp_A_neg_double[0][2] , \out_mux[7][31] , \out_mux[7][30] ,
         \out_mux[7][29] , \out_mux[7][28] , \out_mux[7][27] ,
         \out_mux[7][26] , \out_mux[7][25] , \out_mux[7][24] ,
         \out_mux[7][23] , \out_mux[7][22] , \out_mux[7][21] ,
         \out_mux[7][20] , \out_mux[7][19] , \out_mux[7][18] ,
         \out_mux[7][17] , \out_mux[7][16] , \out_mux[7][15] ,
         \out_mux[7][14] , \out_mux[7][13] , \out_mux[7][12] ,
         \out_mux[7][11] , \out_mux[7][10] , \out_mux[7][9] , \out_mux[7][8] ,
         \out_mux[7][7] , \out_mux[7][6] , \out_mux[7][5] , \out_mux[7][4] ,
         \out_mux[7][3] , \out_mux[7][2] , \out_mux[7][1] , \out_mux[7][0] ,
         \out_mux[6][31] , \out_mux[6][30] , \out_mux[6][29] ,
         \out_mux[6][28] , \out_mux[6][27] , \out_mux[6][26] ,
         \out_mux[6][25] , \out_mux[6][24] , \out_mux[6][23] ,
         \out_mux[6][22] , \out_mux[6][21] , \out_mux[6][20] ,
         \out_mux[6][19] , \out_mux[6][18] , \out_mux[6][17] ,
         \out_mux[6][16] , \out_mux[6][15] , \out_mux[6][14] ,
         \out_mux[6][13] , \out_mux[6][12] , \out_mux[6][11] ,
         \out_mux[6][10] , \out_mux[6][9] , \out_mux[6][8] , \out_mux[6][7] ,
         \out_mux[6][6] , \out_mux[6][5] , \out_mux[6][4] , \out_mux[6][3] ,
         \out_mux[6][2] , \out_mux[6][1] , \out_mux[6][0] , \out_mux[5][31] ,
         \out_mux[5][30] , \out_mux[5][29] , \out_mux[5][28] ,
         \out_mux[5][27] , \out_mux[5][26] , \out_mux[5][25] ,
         \out_mux[5][24] , \out_mux[5][23] , \out_mux[5][22] ,
         \out_mux[5][21] , \out_mux[5][20] , \out_mux[5][19] ,
         \out_mux[5][18] , \out_mux[5][17] , \out_mux[5][16] ,
         \out_mux[5][15] , \out_mux[5][14] , \out_mux[5][13] ,
         \out_mux[5][12] , \out_mux[5][11] , \out_mux[5][10] , \out_mux[5][9] ,
         \out_mux[5][8] , \out_mux[5][7] , \out_mux[5][6] , \out_mux[5][5] ,
         \out_mux[5][4] , \out_mux[5][3] , \out_mux[5][2] , \out_mux[5][1] ,
         \out_mux[5][0] , \out_mux[4][31] , \out_mux[4][30] , \out_mux[4][29] ,
         \out_mux[4][28] , \out_mux[4][27] , \out_mux[4][26] ,
         \out_mux[4][25] , \out_mux[4][24] , \out_mux[4][23] ,
         \out_mux[4][22] , \out_mux[4][21] , \out_mux[4][20] ,
         \out_mux[4][19] , \out_mux[4][18] , \out_mux[4][17] ,
         \out_mux[4][16] , \out_mux[4][15] , \out_mux[4][14] ,
         \out_mux[4][13] , \out_mux[4][12] , \out_mux[4][11] ,
         \out_mux[4][10] , \out_mux[4][9] , \out_mux[4][8] , \out_mux[4][7] ,
         \out_mux[4][6] , \out_mux[4][5] , \out_mux[4][4] , \out_mux[4][3] ,
         \out_mux[4][2] , \out_mux[4][1] , \out_mux[4][0] , \out_mux[3][31] ,
         \out_mux[3][30] , \out_mux[3][29] , \out_mux[3][28] ,
         \out_mux[3][27] , \out_mux[3][26] , \out_mux[3][25] ,
         \out_mux[3][24] , \out_mux[3][23] , \out_mux[3][22] ,
         \out_mux[3][21] , \out_mux[3][20] , \out_mux[3][19] ,
         \out_mux[3][18] , \out_mux[3][17] , \out_mux[3][16] ,
         \out_mux[3][15] , \out_mux[3][14] , \out_mux[3][13] ,
         \out_mux[3][12] , \out_mux[3][11] , \out_mux[3][10] , \out_mux[3][9] ,
         \out_mux[3][8] , \out_mux[3][7] , \out_mux[3][6] , \out_mux[3][5] ,
         \out_mux[3][4] , \out_mux[3][3] , \out_mux[3][2] , \out_mux[3][1] ,
         \out_mux[3][0] , \out_mux[2][31] , \out_mux[2][30] , \out_mux[2][29] ,
         \out_mux[2][28] , \out_mux[2][27] , \out_mux[2][26] ,
         \out_mux[2][25] , \out_mux[2][24] , \out_mux[2][23] ,
         \out_mux[2][22] , \out_mux[2][21] , \out_mux[2][20] ,
         \out_mux[2][19] , \out_mux[2][18] , \out_mux[2][17] ,
         \out_mux[2][16] , \out_mux[2][15] , \out_mux[2][14] ,
         \out_mux[2][13] , \out_mux[2][12] , \out_mux[2][11] ,
         \out_mux[2][10] , \out_mux[2][9] , \out_mux[2][8] , \out_mux[2][7] ,
         \out_mux[2][6] , \out_mux[2][5] , \out_mux[2][4] , \out_mux[2][3] ,
         \out_mux[2][2] , \out_mux[2][1] , \out_mux[2][0] , \out_mux[1][31] ,
         \out_mux[1][30] , \out_mux[1][29] , \out_mux[1][28] ,
         \out_mux[1][27] , \out_mux[1][26] , \out_mux[1][25] ,
         \out_mux[1][24] , \out_mux[1][23] , \out_mux[1][22] ,
         \out_mux[1][21] , \out_mux[1][20] , \out_mux[1][19] ,
         \out_mux[1][18] , \out_mux[1][17] , \out_mux[1][16] ,
         \out_mux[1][15] , \out_mux[1][14] , \out_mux[1][13] ,
         \out_mux[1][12] , \out_mux[1][11] , \out_mux[1][10] , \out_mux[1][9] ,
         \out_mux[1][8] , \out_mux[1][7] , \out_mux[1][6] , \out_mux[1][5] ,
         \out_mux[1][4] , \out_mux[1][3] , \out_mux[1][2] , \out_mux[1][1] ,
         \out_mux[1][0] , \out_mux[0][31] , \out_mux[0][30] , \out_mux[0][29] ,
         \out_mux[0][28] , \out_mux[0][27] , \out_mux[0][26] ,
         \out_mux[0][25] , \out_mux[0][24] , \out_mux[0][23] ,
         \out_mux[0][22] , \out_mux[0][21] , \out_mux[0][20] ,
         \out_mux[0][19] , \out_mux[0][18] , \out_mux[0][17] ,
         \out_mux[0][16] , \out_mux[0][15] , \out_mux[0][14] ,
         \out_mux[0][13] , \out_mux[0][12] , \out_mux[0][11] ,
         \out_mux[0][10] , \out_mux[0][9] , \out_mux[0][8] , \out_mux[0][7] ,
         \out_mux[0][6] , \out_mux[0][5] , \out_mux[0][4] , \out_mux[0][3] ,
         \out_mux[0][2] , \out_mux[0][1] , \out_mux[0][0] , \out_sum[5][31] ,
         \out_sum[5][30] , \out_sum[5][29] , \out_sum[5][28] ,
         \out_sum[5][27] , \out_sum[5][26] , \out_sum[5][25] ,
         \out_sum[5][24] , \out_sum[5][23] , \out_sum[5][22] ,
         \out_sum[5][21] , \out_sum[5][20] , \out_sum[5][19] ,
         \out_sum[5][18] , \out_sum[5][17] , \out_sum[5][16] ,
         \out_sum[5][15] , \out_sum[5][14] , \out_sum[5][13] ,
         \out_sum[5][12] , \out_sum[5][11] , \out_sum[5][10] , \out_sum[5][9] ,
         \out_sum[5][8] , \out_sum[5][7] , \out_sum[5][6] , \out_sum[5][5] ,
         \out_sum[5][4] , \out_sum[5][3] , \out_sum[5][2] , \out_sum[5][1] ,
         \out_sum[5][0] , \out_sum[4][31] , \out_sum[4][30] , \out_sum[4][29] ,
         \out_sum[4][28] , \out_sum[4][27] , \out_sum[4][26] ,
         \out_sum[4][25] , \out_sum[4][24] , \out_sum[4][23] ,
         \out_sum[4][22] , \out_sum[4][21] , \out_sum[4][20] ,
         \out_sum[4][19] , \out_sum[4][18] , \out_sum[4][17] ,
         \out_sum[4][16] , \out_sum[4][15] , \out_sum[4][14] ,
         \out_sum[4][13] , \out_sum[4][12] , \out_sum[4][11] ,
         \out_sum[4][10] , \out_sum[4][9] , \out_sum[4][8] , \out_sum[4][7] ,
         \out_sum[4][6] , \out_sum[4][5] , \out_sum[4][4] , \out_sum[4][3] ,
         \out_sum[4][2] , \out_sum[4][1] , \out_sum[4][0] , \out_sum[3][31] ,
         \out_sum[3][30] , \out_sum[3][29] , \out_sum[3][28] ,
         \out_sum[3][27] , \out_sum[3][26] , \out_sum[3][25] ,
         \out_sum[3][24] , \out_sum[3][23] , \out_sum[3][22] ,
         \out_sum[3][21] , \out_sum[3][20] , \out_sum[3][19] ,
         \out_sum[3][18] , \out_sum[3][17] , \out_sum[3][16] ,
         \out_sum[3][15] , \out_sum[3][14] , \out_sum[3][13] ,
         \out_sum[3][12] , \out_sum[3][11] , \out_sum[3][10] , \out_sum[3][9] ,
         \out_sum[3][8] , \out_sum[3][7] , \out_sum[3][6] , \out_sum[3][5] ,
         \out_sum[3][4] , \out_sum[3][3] , \out_sum[3][2] , \out_sum[3][1] ,
         \out_sum[3][0] , \out_sum[2][31] , \out_sum[2][30] , \out_sum[2][29] ,
         \out_sum[2][28] , \out_sum[2][27] , \out_sum[2][26] ,
         \out_sum[2][25] , \out_sum[2][24] , \out_sum[2][23] ,
         \out_sum[2][22] , \out_sum[2][21] , \out_sum[2][20] ,
         \out_sum[2][19] , \out_sum[2][18] , \out_sum[2][17] ,
         \out_sum[2][16] , \out_sum[2][15] , \out_sum[2][14] ,
         \out_sum[2][13] , \out_sum[2][12] , \out_sum[2][11] ,
         \out_sum[2][10] , \out_sum[2][9] , \out_sum[2][8] , \out_sum[2][7] ,
         \out_sum[2][6] , \out_sum[2][5] , \out_sum[2][4] , \out_sum[2][3] ,
         \out_sum[2][2] , \out_sum[2][1] , \out_sum[2][0] , \out_sum[1][31] ,
         \out_sum[1][30] , \out_sum[1][29] , \out_sum[1][28] ,
         \out_sum[1][27] , \out_sum[1][26] , \out_sum[1][25] ,
         \out_sum[1][24] , \out_sum[1][23] , \out_sum[1][22] ,
         \out_sum[1][21] , \out_sum[1][20] , \out_sum[1][19] ,
         \out_sum[1][18] , \out_sum[1][17] , \out_sum[1][16] ,
         \out_sum[1][15] , \out_sum[1][14] , \out_sum[1][13] ,
         \out_sum[1][12] , \out_sum[1][11] , \out_sum[1][10] , \out_sum[1][9] ,
         \out_sum[1][8] , \out_sum[1][7] , \out_sum[1][6] , \out_sum[1][5] ,
         \out_sum[1][4] , \out_sum[1][3] , \out_sum[1][2] , \out_sum[1][1] ,
         \out_sum[1][0] , \out_sum[0][31] , \out_sum[0][30] , \out_sum[0][29] ,
         \out_sum[0][28] , \out_sum[0][27] , \out_sum[0][26] ,
         \out_sum[0][25] , \out_sum[0][24] , \out_sum[0][23] ,
         \out_sum[0][22] , \out_sum[0][21] , \out_sum[0][20] ,
         \out_sum[0][19] , \out_sum[0][18] , \out_sum[0][17] ,
         \out_sum[0][16] , \out_sum[0][15] , \out_sum[0][14] ,
         \out_sum[0][13] , \out_sum[0][12] , \out_sum[0][11] ,
         \out_sum[0][10] , \out_sum[0][9] , \out_sum[0][8] , \out_sum[0][7] ,
         \out_sum[0][6] , \out_sum[0][5] , \out_sum[0][4] , \out_sum[0][3] ,
         \out_sum[0][2] , \out_sum[0][1] , \out_sum[0][0] ,
         \add_83_2_C132_G8/carry[17] , \add_83_2_C132_G8/carry[18] ,
         \add_83_2_C132_G8/carry[19] , \add_83_2_C132_G8/carry[20] ,
         \add_83_2_C132_G8/carry[21] , \add_83_2_C132_G8/carry[22] ,
         \add_83_2_C132_G8/carry[23] , \add_83_2_C132_G8/carry[24] ,
         \add_83_2_C132_G8/carry[25] , \add_83_2_C132_G8/carry[26] ,
         \add_83_2_C132_G8/carry[27] , \add_83_2_C132_G8/carry[28] ,
         \add_83_2_C132_G8/carry[29] , \add_83_2_C132_G8/carry[30] ,
         \add_83_2_C132_G8/carry[31] , \add_83_2_C130_G8/carry[15] ,
         \add_83_2_C130_G8/carry[16] , \add_83_2_C130_G8/carry[17] ,
         \add_83_2_C130_G8/carry[18] , \add_83_2_C130_G8/carry[19] ,
         \add_83_2_C130_G8/carry[20] , \add_83_2_C130_G8/carry[21] ,
         \add_83_2_C130_G8/carry[22] , \add_83_2_C130_G8/carry[23] ,
         \add_83_2_C130_G8/carry[24] , \add_83_2_C130_G8/carry[25] ,
         \add_83_2_C130_G8/carry[26] , \add_83_2_C130_G8/carry[27] ,
         \add_83_2_C130_G8/carry[28] , \add_83_2_C130_G8/carry[29] ,
         \add_83_2_C130_G8/carry[30] , \add_83_2_C130_G8/carry[31] ,
         \add_83_2_C132_G7/carry[15] , \add_83_2_C132_G7/carry[16] ,
         \add_83_2_C132_G7/carry[17] , \add_83_2_C132_G7/carry[18] ,
         \add_83_2_C132_G7/carry[19] , \add_83_2_C132_G7/carry[20] ,
         \add_83_2_C132_G7/carry[21] , \add_83_2_C132_G7/carry[22] ,
         \add_83_2_C132_G7/carry[23] , \add_83_2_C132_G7/carry[24] ,
         \add_83_2_C132_G7/carry[25] , \add_83_2_C132_G7/carry[26] ,
         \add_83_2_C132_G7/carry[27] , \add_83_2_C132_G7/carry[28] ,
         \add_83_2_C132_G7/carry[29] , \add_83_2_C132_G7/carry[30] ,
         \add_83_2_C132_G7/carry[31] , \add_83_2_C130_G7/carry[14] ,
         \add_83_2_C130_G7/carry[15] , \add_83_2_C130_G7/carry[16] ,
         \add_83_2_C130_G7/carry[17] , \add_83_2_C130_G7/carry[18] ,
         \add_83_2_C130_G7/carry[19] , \add_83_2_C130_G7/carry[20] ,
         \add_83_2_C130_G7/carry[21] , \add_83_2_C130_G7/carry[22] ,
         \add_83_2_C130_G7/carry[23] , \add_83_2_C130_G7/carry[24] ,
         \add_83_2_C130_G7/carry[25] , \add_83_2_C130_G7/carry[26] ,
         \add_83_2_C130_G7/carry[27] , \add_83_2_C130_G7/carry[28] ,
         \add_83_2_C130_G7/carry[29] , \add_83_2_C130_G7/carry[30] ,
         \add_83_2_C130_G7/carry[31] , \add_83_2_C132_G5/carry[11] ,
         \add_83_2_C132_G5/carry[12] , \add_83_2_C132_G5/carry[13] ,
         \add_83_2_C132_G5/carry[14] , \add_83_2_C132_G5/carry[15] ,
         \add_83_2_C132_G5/carry[16] , \add_83_2_C132_G5/carry[17] ,
         \add_83_2_C132_G5/carry[18] , \add_83_2_C132_G5/carry[19] ,
         \add_83_2_C132_G5/carry[20] , \add_83_2_C132_G5/carry[21] ,
         \add_83_2_C132_G5/carry[22] , \add_83_2_C132_G5/carry[23] ,
         \add_83_2_C132_G5/carry[24] , \add_83_2_C130_G5/carry[10] ,
         \add_83_2_C130_G5/carry[11] , \add_83_2_C130_G5/carry[12] ,
         \add_83_2_C130_G5/carry[13] , \add_83_2_C130_G5/carry[14] ,
         \add_83_2_C130_G5/carry[15] , \add_83_2_C130_G5/carry[16] ,
         \add_83_2_C130_G5/carry[17] , \add_83_2_C130_G5/carry[18] ,
         \add_83_2_C130_G5/carry[19] , \add_83_2_C130_G5/carry[20] ,
         \add_83_2_C130_G5/carry[21] , \add_83_2_C130_G5/carry[22] ,
         \add_83_2_C130_G5/carry[23] , \add_83_2_C132_G4/carry[9] ,
         \add_83_2_C132_G4/carry[10] , \add_83_2_C132_G4/carry[11] ,
         \add_83_2_C132_G4/carry[12] , \add_83_2_C132_G4/carry[13] ,
         \add_83_2_C132_G4/carry[14] , \add_83_2_C132_G4/carry[15] ,
         \add_83_2_C132_G4/carry[16] , \add_83_2_C132_G4/carry[17] ,
         \add_83_2_C132_G4/carry[18] , \add_83_2_C132_G4/carry[19] ,
         \add_83_2_C132_G4/carry[20] , \add_83_2_C132_G4/carry[21] ,
         \add_83_2_C132_G4/carry[22] , \add_83_2_C130_G4/carry[8] ,
         \add_83_2_C130_G4/carry[9] , \add_83_2_C130_G4/carry[10] ,
         \add_83_2_C130_G4/carry[11] , \add_83_2_C130_G4/carry[12] ,
         \add_83_2_C130_G4/carry[13] , \add_83_2_C130_G4/carry[14] ,
         \add_83_2_C130_G4/carry[15] , \add_83_2_C130_G4/carry[16] ,
         \add_83_2_C130_G4/carry[17] , \add_83_2_C130_G4/carry[18] ,
         \add_83_2_C130_G4/carry[19] , \add_83_2_C130_G4/carry[20] ,
         \add_83_2_C130_G4/carry[21] , \add_83_2_C132_G3/carry[7] ,
         \add_83_2_C132_G3/carry[8] , \add_83_2_C132_G3/carry[9] ,
         \add_83_2_C132_G3/carry[10] , \add_83_2_C132_G3/carry[11] ,
         \add_83_2_C132_G3/carry[12] , \add_83_2_C132_G3/carry[13] ,
         \add_83_2_C132_G3/carry[14] , \add_83_2_C132_G3/carry[15] ,
         \add_83_2_C132_G3/carry[16] , \add_83_2_C132_G3/carry[17] ,
         \add_83_2_C132_G3/carry[18] , \add_83_2_C132_G3/carry[19] ,
         \add_83_2_C132_G3/carry[20] , \add_83_2_C130_G3/carry[6] ,
         \add_83_2_C130_G3/carry[7] , \add_83_2_C130_G3/carry[8] ,
         \add_83_2_C130_G3/carry[9] , \add_83_2_C130_G3/carry[10] ,
         \add_83_2_C130_G3/carry[11] , \add_83_2_C130_G3/carry[12] ,
         \add_83_2_C130_G3/carry[13] , \add_83_2_C130_G3/carry[14] ,
         \add_83_2_C130_G3/carry[15] , \add_83_2_C130_G3/carry[16] ,
         \add_83_2_C130_G3/carry[17] , \add_83_2_C130_G3/carry[18] ,
         \add_83_2_C130_G3/carry[19] , \add_83_2_C132_G2/carry[5] ,
         \add_83_2_C132_G2/carry[6] , \add_83_2_C132_G2/carry[7] ,
         \add_83_2_C132_G2/carry[8] , \add_83_2_C132_G2/carry[9] ,
         \add_83_2_C132_G2/carry[10] , \add_83_2_C132_G2/carry[11] ,
         \add_83_2_C132_G2/carry[12] , \add_83_2_C132_G2/carry[13] ,
         \add_83_2_C132_G2/carry[16] , \add_83_2_C132_G2/carry[17] ,
         \add_83_2_C132_G2/carry[18] , \add_83_2_C130_G2/carry[4] ,
         \add_83_2_C130_G2/carry[5] , \add_83_2_C130_G2/carry[6] ,
         \add_83_2_C130_G2/carry[7] , \add_83_2_C130_G2/carry[8] ,
         \add_83_2_C130_G2/carry[9] , \add_83_2_C130_G2/carry[10] ,
         \add_83_2_C130_G2/carry[11] , \add_83_2_C130_G2/carry[12] ,
         \add_83_2_C130_G2/carry[13] , \add_83_2_C130_G2/carry[14] ,
         \add_83_2_C130_G2/carry[15] , \add_83_2_C130_G2/carry[16] ,
         \add_83_2_C130_G2/carry[17] , \add_83_2_C111/carry[6] ,
         \add_83_2_C111/carry[7] , \add_83_2_C111/carry[10] ,
         \add_83_2_C111/carry[16] , \add_109/carry[2] , \add_109/carry[4] ,
         \add_109/carry[5] , \add_109/carry[6] , \add_109/carry[8] ,
         \add_109/carry[12] , \add_109/carry[15] , n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20;

  booth_mux_generic_N32_0 Muxes_0 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n69, n69, n69, n69, n69, n69, n69, n69, n69, n68, 
        n68, n68, n68, n68, n68, n68, n68, A[14:0]}), .A_neg({n52, n52, n52, 
        n52, n52, n52, n52, n52, n52, n52, n52, \tmp_A_neg[0][31] , n52, n52, 
        \tmp_A_neg[0][31] , \tmp_A_neg[0][31] , \tmp_A_neg[0][15] , 
        \tmp_A_neg[0][14] , \tmp_A_neg[0][13] , \tmp_A_neg[0][12] , 
        \tmp_A_neg[0][11] , \tmp_A_neg[0][10] , \tmp_A_neg[0][9] , 
        \tmp_A_neg[0][8] , \tmp_A_neg[0][7] , \tmp_A_neg[0][6] , 
        \tmp_A_neg[0][5] , \tmp_A_neg[0][4] , \tmp_A_neg[0][3] , 
        \tmp_A_neg[0][2] , \tmp_A_neg[0][1] , A[0]}), .A_double({n68, n68, n68, 
        n68, n68, n67, n67, n67, n67, n67, n67, n67, n67, n67, n67, n67, 
        A[14:1], n55, 1'b0}), .A_neg_double({\tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][31] , \tmp_A_neg_double[0][31] , 
        \tmp_A_neg_double[0][16] , \tmp_A_neg_double[0][15] , 
        \tmp_A_neg_double[0][14] , \tmp_A_neg_double[0][13] , 
        \tmp_A_neg_double[0][12] , \tmp_A_neg_double[0][11] , 
        \tmp_A_neg_double[0][10] , \tmp_A_neg_double[0][9] , 
        \tmp_A_neg_double[0][8] , \tmp_A_neg_double[0][7] , 
        \tmp_A_neg_double[0][6] , \tmp_A_neg_double[0][5] , 
        \tmp_A_neg_double[0][4] , \tmp_A_neg_double[0][3] , 
        \tmp_A_neg_double[0][2] , n55, 1'b0}), .SEL({B[1:0], 1'b0}), .Y({
        \out_mux[0][31] , \out_mux[0][30] , \out_mux[0][29] , \out_mux[0][28] , 
        \out_mux[0][27] , \out_mux[0][26] , \out_mux[0][25] , \out_mux[0][24] , 
        \out_mux[0][23] , \out_mux[0][22] , \out_mux[0][21] , \out_mux[0][20] , 
        \out_mux[0][19] , \out_mux[0][18] , \out_mux[0][17] , \out_mux[0][16] , 
        \out_mux[0][15] , \out_mux[0][14] , \out_mux[0][13] , \out_mux[0][12] , 
        \out_mux[0][11] , \out_mux[0][10] , \out_mux[0][9] , \out_mux[0][8] , 
        \out_mux[0][7] , \out_mux[0][6] , \out_mux[0][5] , \out_mux[0][4] , 
        \out_mux[0][3] , \out_mux[0][2] , \out_mux[0][1] , \out_mux[0][0] })
         );
  booth_mux_generic_N32_7 Muxes_1 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n60, n60, n60, n59, n59, n59, n59, n59, n59, n59, 
        n59, n59, n59, n59, n59, A[14:1], n55, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , 
        \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , 
        \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , 
        \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , 
        \tmp_A_neg[1][31] , \tmp_A_neg[1][31] , \tmp_A_neg[1][17] , 
        \tmp_A_neg[1][16] , \tmp_A_neg[1][15] , \tmp_A_neg[1][14] , 
        \tmp_A_neg[1][13] , \tmp_A_neg[1][12] , \tmp_A_neg[1][11] , 
        \tmp_A_neg[1][10] , \tmp_A_neg[1][9] , \tmp_A_neg[1][8] , 
        \tmp_A_neg[1][7] , \tmp_A_neg[1][6] , \tmp_A_neg[1][5] , 
        \tmp_A_neg[1][4] , \tmp_A_neg[1][3] , n55, 1'b0, 1'b0}), .A_double({
        n59, n58, n58, n58, n58, n58, n58, n58, n58, n58, n58, n58, n58, n58, 
        A[14:1], n55, 1'b0, 1'b0, 1'b0}), .A_neg_double({n45, n45, n45, n45, 
        n45, n45, n45, n45, n45, n45, n45, n45, \tmp_A_neg_double[1][31] , 
        \tmp_A_neg_double[1][18] , \tmp_A_neg_double[1][17] , 
        \tmp_A_neg_double[1][16] , \tmp_A_neg_double[1][15] , 
        \tmp_A_neg_double[1][14] , \tmp_A_neg_double[1][13] , 
        \tmp_A_neg_double[1][12] , \tmp_A_neg_double[1][11] , 
        \tmp_A_neg_double[1][10] , \tmp_A_neg_double[1][9] , 
        \tmp_A_neg_double[1][8] , \tmp_A_neg_double[1][7] , 
        \tmp_A_neg_double[1][6] , \tmp_A_neg_double[1][5] , 
        \tmp_A_neg_double[1][4] , n55, 1'b0, 1'b0, 1'b0}), .SEL(B[3:1]), .Y({
        \out_mux[1][31] , \out_mux[1][30] , \out_mux[1][29] , \out_mux[1][28] , 
        \out_mux[1][27] , \out_mux[1][26] , \out_mux[1][25] , \out_mux[1][24] , 
        \out_mux[1][23] , \out_mux[1][22] , \out_mux[1][21] , \out_mux[1][20] , 
        \out_mux[1][19] , \out_mux[1][18] , \out_mux[1][17] , \out_mux[1][16] , 
        \out_mux[1][15] , \out_mux[1][14] , \out_mux[1][13] , \out_mux[1][12] , 
        \out_mux[1][11] , \out_mux[1][10] , \out_mux[1][9] , \out_mux[1][8] , 
        \out_mux[1][7] , \out_mux[1][6] , \out_mux[1][5] , \out_mux[1][4] , 
        \out_mux[1][3] , \out_mux[1][2] , \out_mux[1][1] , \out_mux[1][0] })
         );
  P4adder_N32_PowerN5_0 sum_1 ( .A({\out_mux[1][31] , \out_mux[1][30] , 
        \out_mux[1][29] , \out_mux[1][28] , \out_mux[1][27] , \out_mux[1][26] , 
        \out_mux[1][25] , \out_mux[1][24] , \out_mux[1][23] , \out_mux[1][22] , 
        \out_mux[1][21] , \out_mux[1][20] , \out_mux[1][19] , \out_mux[1][18] , 
        \out_mux[1][17] , \out_mux[1][16] , \out_mux[1][15] , \out_mux[1][14] , 
        \out_mux[1][13] , \out_mux[1][12] , \out_mux[1][11] , \out_mux[1][10] , 
        \out_mux[1][9] , \out_mux[1][8] , \out_mux[1][7] , \out_mux[1][6] , 
        \out_mux[1][5] , \out_mux[1][4] , \out_mux[1][3] , \out_mux[1][2] , 
        \out_mux[1][1] , \out_mux[1][0] }), .B({\out_mux[0][31] , 
        \out_mux[0][30] , \out_mux[0][29] , \out_mux[0][28] , \out_mux[0][27] , 
        \out_mux[0][26] , \out_mux[0][25] , \out_mux[0][24] , \out_mux[0][23] , 
        \out_mux[0][22] , \out_mux[0][21] , \out_mux[0][20] , \out_mux[0][19] , 
        \out_mux[0][18] , \out_mux[0][17] , \out_mux[0][16] , \out_mux[0][15] , 
        \out_mux[0][14] , \out_mux[0][13] , \out_mux[0][12] , \out_mux[0][11] , 
        \out_mux[0][10] , \out_mux[0][9] , \out_mux[0][8] , \out_mux[0][7] , 
        \out_mux[0][6] , \out_mux[0][5] , \out_mux[0][4] , \out_mux[0][3] , 
        \out_mux[0][2] , \out_mux[0][1] , \out_mux[0][0] }), .Ci(1'b0), .S({
        \out_sum[0][31] , \out_sum[0][30] , \out_sum[0][29] , \out_sum[0][28] , 
        \out_sum[0][27] , \out_sum[0][26] , \out_sum[0][25] , \out_sum[0][24] , 
        \out_sum[0][23] , \out_sum[0][22] , \out_sum[0][21] , \out_sum[0][20] , 
        \out_sum[0][19] , \out_sum[0][18] , \out_sum[0][17] , \out_sum[0][16] , 
        \out_sum[0][15] , \out_sum[0][14] , \out_sum[0][13] , \out_sum[0][12] , 
        \out_sum[0][11] , \out_sum[0][10] , \out_sum[0][9] , \out_sum[0][8] , 
        \out_sum[0][7] , \out_sum[0][6] , \out_sum[0][5] , \out_sum[0][4] , 
        \out_sum[0][3] , \out_sum[0][2] , \out_sum[0][1] , \out_sum[0][0] })
         );
  booth_mux_generic_N32_6 Muxes_2 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n62, n62, n61, n61, n61, n61, n61, n61, n61, n61, 
        n61, n61, n61, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , 
        \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , 
        \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , 
        \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , \tmp_A_neg[2][31] , 
        \tmp_A_neg[2][19] , \tmp_A_neg[2][18] , \tmp_A_neg[2][17] , 
        \tmp_A_neg[2][16] , \tmp_A_neg[2][15] , \tmp_A_neg[2][14] , 
        \tmp_A_neg[2][13] , \tmp_A_neg[2][12] , \tmp_A_neg[2][11] , 
        \tmp_A_neg[2][10] , \tmp_A_neg[2][9] , \tmp_A_neg[2][8] , 
        \tmp_A_neg[2][7] , \tmp_A_neg[2][6] , \tmp_A_neg[2][5] , A[0], 1'b0, 
        1'b0, 1'b0, 1'b0}), .A_double({n61, n61, n60, n60, n60, n60, n60, n60, 
        n60, n60, n60, n60, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .A_neg_double({\tmp_A_neg_double[2][31] , \tmp_A_neg_double[2][31] , 
        \tmp_A_neg_double[2][31] , \tmp_A_neg_double[2][31] , 
        \tmp_A_neg_double[2][31] , \tmp_A_neg_double[2][31] , 
        \tmp_A_neg_double[2][31] , \tmp_A_neg_double[2][31] , 
        \tmp_A_neg_double[2][31] , \tmp_A_neg_double[2][31] , 
        \tmp_A_neg_double[2][31] , \tmp_A_neg_double[2][20] , 
        \tmp_A_neg_double[2][19] , \tmp_A_neg_double[2][18] , 
        \tmp_A_neg_double[2][17] , \tmp_A_neg_double[2][16] , 
        \tmp_A_neg_double[2][15] , \tmp_A_neg_double[2][14] , 
        \tmp_A_neg_double[2][13] , \tmp_A_neg_double[2][12] , 
        \tmp_A_neg_double[2][11] , \tmp_A_neg_double[2][10] , 
        \tmp_A_neg_double[2][9] , \tmp_A_neg_double[2][8] , 
        \tmp_A_neg_double[2][7] , \tmp_A_neg_double[2][6] , A[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(B[5:3]), .Y({\out_mux[2][31] , 
        \out_mux[2][30] , \out_mux[2][29] , \out_mux[2][28] , \out_mux[2][27] , 
        \out_mux[2][26] , \out_mux[2][25] , \out_mux[2][24] , \out_mux[2][23] , 
        \out_mux[2][22] , \out_mux[2][21] , \out_mux[2][20] , \out_mux[2][19] , 
        \out_mux[2][18] , \out_mux[2][17] , \out_mux[2][16] , \out_mux[2][15] , 
        \out_mux[2][14] , \out_mux[2][13] , \out_mux[2][12] , \out_mux[2][11] , 
        \out_mux[2][10] , \out_mux[2][9] , \out_mux[2][8] , \out_mux[2][7] , 
        \out_mux[2][6] , \out_mux[2][5] , \out_mux[2][4] , \out_mux[2][3] , 
        \out_mux[2][2] , \out_mux[2][1] , \out_mux[2][0] }) );
  P4adder_N32_PowerN5_6 sum_2 ( .A({\out_mux[2][31] , \out_mux[2][30] , 
        \out_mux[2][29] , \out_mux[2][28] , \out_mux[2][27] , \out_mux[2][26] , 
        \out_mux[2][25] , \out_mux[2][24] , \out_mux[2][23] , \out_mux[2][22] , 
        \out_mux[2][21] , \out_mux[2][20] , \out_mux[2][19] , \out_mux[2][18] , 
        \out_mux[2][17] , \out_mux[2][16] , \out_mux[2][15] , \out_mux[2][14] , 
        \out_mux[2][13] , \out_mux[2][12] , \out_mux[2][11] , \out_mux[2][10] , 
        \out_mux[2][9] , \out_mux[2][8] , \out_mux[2][7] , \out_mux[2][6] , 
        \out_mux[2][5] , \out_mux[2][4] , \out_mux[2][3] , \out_mux[2][2] , 
        \out_mux[2][1] , \out_mux[2][0] }), .B({\out_sum[0][31] , 
        \out_sum[0][30] , \out_sum[0][29] , \out_sum[0][28] , \out_sum[0][27] , 
        \out_sum[0][26] , \out_sum[0][25] , \out_sum[0][24] , \out_sum[0][23] , 
        \out_sum[0][22] , \out_sum[0][21] , \out_sum[0][20] , \out_sum[0][19] , 
        \out_sum[0][18] , \out_sum[0][17] , \out_sum[0][16] , \out_sum[0][15] , 
        \out_sum[0][14] , \out_sum[0][13] , \out_sum[0][12] , \out_sum[0][11] , 
        \out_sum[0][10] , \out_sum[0][9] , \out_sum[0][8] , \out_sum[0][7] , 
        \out_sum[0][6] , \out_sum[0][5] , \out_sum[0][4] , \out_sum[0][3] , 
        \out_sum[0][2] , \out_sum[0][1] , \out_sum[0][0] }), .Ci(1'b0), .S({
        \out_sum[1][31] , \out_sum[1][30] , \out_sum[1][29] , \out_sum[1][28] , 
        \out_sum[1][27] , \out_sum[1][26] , \out_sum[1][25] , \out_sum[1][24] , 
        \out_sum[1][23] , \out_sum[1][22] , \out_sum[1][21] , \out_sum[1][20] , 
        \out_sum[1][19] , \out_sum[1][18] , \out_sum[1][17] , \out_sum[1][16] , 
        \out_sum[1][15] , \out_sum[1][14] , \out_sum[1][13] , \out_sum[1][12] , 
        \out_sum[1][11] , \out_sum[1][10] , \out_sum[1][9] , \out_sum[1][8] , 
        \out_sum[1][7] , \out_sum[1][6] , \out_sum[1][5] , \out_sum[1][4] , 
        \out_sum[1][3] , \out_sum[1][2] , \out_sum[1][1] , \out_sum[1][0] })
         );
  booth_mux_generic_N32_5 Muxes_3 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n63, n63, n63, n63, n63, n63, n63, n63, n63, n63, 
        n62, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[3][31] , \tmp_A_neg[3][31] , \tmp_A_neg[3][31] , 
        \tmp_A_neg[3][31] , \tmp_A_neg[3][31] , \tmp_A_neg[3][31] , 
        \tmp_A_neg[3][31] , \tmp_A_neg[3][31] , \tmp_A_neg[3][31] , 
        \tmp_A_neg[3][31] , \tmp_A_neg[3][21] , \tmp_A_neg[3][20] , 
        \tmp_A_neg[3][19] , \tmp_A_neg[3][18] , \tmp_A_neg[3][17] , 
        \tmp_A_neg[3][16] , \tmp_A_neg[3][15] , \tmp_A_neg[3][14] , 
        \tmp_A_neg[3][13] , \tmp_A_neg[3][12] , \tmp_A_neg[3][11] , 
        \tmp_A_neg[3][10] , \tmp_A_neg[3][9] , \tmp_A_neg[3][8] , 
        \tmp_A_neg[3][7] , A[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .A_double({n62, n62, n62, n62, n62, n62, n62, n62, n62, n62, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg_double({
        \tmp_A_neg_double[3][31] , \tmp_A_neg_double[3][31] , 
        \tmp_A_neg_double[3][31] , \tmp_A_neg_double[3][31] , 
        \tmp_A_neg_double[3][31] , \tmp_A_neg_double[3][31] , 
        \tmp_A_neg_double[3][31] , \tmp_A_neg_double[3][31] , 
        \tmp_A_neg_double[3][31] , \tmp_A_neg_double[3][22] , 
        \tmp_A_neg_double[3][21] , \tmp_A_neg_double[3][20] , 
        \tmp_A_neg_double[3][19] , \tmp_A_neg_double[3][18] , 
        \tmp_A_neg_double[3][17] , \tmp_A_neg_double[3][16] , 
        \tmp_A_neg_double[3][15] , \tmp_A_neg_double[3][14] , 
        \tmp_A_neg_double[3][13] , \tmp_A_neg_double[3][12] , 
        \tmp_A_neg_double[3][11] , \tmp_A_neg_double[3][10] , 
        \tmp_A_neg_double[3][9] , \tmp_A_neg_double[3][8] , A[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(B[7:5]), .Y({\out_mux[3][31] , 
        \out_mux[3][30] , \out_mux[3][29] , \out_mux[3][28] , \out_mux[3][27] , 
        \out_mux[3][26] , \out_mux[3][25] , \out_mux[3][24] , \out_mux[3][23] , 
        \out_mux[3][22] , \out_mux[3][21] , \out_mux[3][20] , \out_mux[3][19] , 
        \out_mux[3][18] , \out_mux[3][17] , \out_mux[3][16] , \out_mux[3][15] , 
        \out_mux[3][14] , \out_mux[3][13] , \out_mux[3][12] , \out_mux[3][11] , 
        \out_mux[3][10] , \out_mux[3][9] , \out_mux[3][8] , \out_mux[3][7] , 
        \out_mux[3][6] , \out_mux[3][5] , \out_mux[3][4] , \out_mux[3][3] , 
        \out_mux[3][2] , \out_mux[3][1] , \out_mux[3][0] }) );
  P4adder_N32_PowerN5_5 sum_3 ( .A({\out_mux[3][31] , \out_mux[3][30] , 
        \out_mux[3][29] , \out_mux[3][28] , \out_mux[3][27] , \out_mux[3][26] , 
        \out_mux[3][25] , \out_mux[3][24] , \out_mux[3][23] , \out_mux[3][22] , 
        \out_mux[3][21] , \out_mux[3][20] , \out_mux[3][19] , \out_mux[3][18] , 
        \out_mux[3][17] , \out_mux[3][16] , \out_mux[3][15] , \out_mux[3][14] , 
        \out_mux[3][13] , \out_mux[3][12] , \out_mux[3][11] , \out_mux[3][10] , 
        \out_mux[3][9] , \out_mux[3][8] , \out_mux[3][7] , \out_mux[3][6] , 
        \out_mux[3][5] , \out_mux[3][4] , \out_mux[3][3] , \out_mux[3][2] , 
        \out_mux[3][1] , \out_mux[3][0] }), .B({\out_sum[1][31] , 
        \out_sum[1][30] , \out_sum[1][29] , \out_sum[1][28] , \out_sum[1][27] , 
        \out_sum[1][26] , \out_sum[1][25] , \out_sum[1][24] , \out_sum[1][23] , 
        \out_sum[1][22] , \out_sum[1][21] , \out_sum[1][20] , \out_sum[1][19] , 
        \out_sum[1][18] , \out_sum[1][17] , \out_sum[1][16] , \out_sum[1][15] , 
        \out_sum[1][14] , \out_sum[1][13] , \out_sum[1][12] , \out_sum[1][11] , 
        \out_sum[1][10] , \out_sum[1][9] , \out_sum[1][8] , \out_sum[1][7] , 
        \out_sum[1][6] , \out_sum[1][5] , \out_sum[1][4] , \out_sum[1][3] , 
        \out_sum[1][2] , \out_sum[1][1] , \out_sum[1][0] }), .Ci(1'b0), .S({
        \out_sum[2][31] , \out_sum[2][30] , \out_sum[2][29] , \out_sum[2][28] , 
        \out_sum[2][27] , \out_sum[2][26] , \out_sum[2][25] , \out_sum[2][24] , 
        \out_sum[2][23] , \out_sum[2][22] , \out_sum[2][21] , \out_sum[2][20] , 
        \out_sum[2][19] , \out_sum[2][18] , \out_sum[2][17] , \out_sum[2][16] , 
        \out_sum[2][15] , \out_sum[2][14] , \out_sum[2][13] , \out_sum[2][12] , 
        \out_sum[2][11] , \out_sum[2][10] , \out_sum[2][9] , \out_sum[2][8] , 
        \out_sum[2][7] , \out_sum[2][6] , \out_sum[2][5] , \out_sum[2][4] , 
        \out_sum[2][3] , \out_sum[2][2] , \out_sum[2][1] , \out_sum[2][0] })
         );
  booth_mux_generic_N32_4 Muxes_4 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n65, n64, n64, n64, n64, n64, n64, n64, n64, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[4][31] , \tmp_A_neg[4][31] , \tmp_A_neg[4][31] , 
        \tmp_A_neg[4][31] , \tmp_A_neg[4][31] , \tmp_A_neg[4][31] , 
        \tmp_A_neg[4][31] , \tmp_A_neg[4][31] , \tmp_A_neg[4][23] , 
        \tmp_A_neg[4][22] , \tmp_A_neg[4][21] , \tmp_A_neg[4][20] , 
        \tmp_A_neg[4][19] , \tmp_A_neg[4][18] , \tmp_A_neg[4][17] , 
        \tmp_A_neg[4][16] , \tmp_A_neg[4][15] , \tmp_A_neg[4][14] , 
        \tmp_A_neg[4][13] , \tmp_A_neg[4][12] , \tmp_A_neg[4][11] , 
        \tmp_A_neg[4][10] , \tmp_A_neg[4][9] , A[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_double({n64, n64, n64, n64, n64, n63, n63, 
        n63, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .A_neg_double({\tmp_A_neg_double[4][31] , \tmp_A_neg_double[4][31] , 
        \tmp_A_neg_double[4][31] , \tmp_A_neg_double[4][31] , 
        \tmp_A_neg_double[4][31] , \tmp_A_neg_double[4][31] , 
        \tmp_A_neg_double[4][31] , \tmp_A_neg_double[4][24] , 
        \tmp_A_neg_double[4][23] , \tmp_A_neg_double[4][22] , 
        \tmp_A_neg_double[4][21] , \tmp_A_neg_double[4][20] , 
        \tmp_A_neg_double[4][19] , \tmp_A_neg_double[4][18] , 
        \tmp_A_neg_double[4][17] , \tmp_A_neg_double[4][16] , 
        \tmp_A_neg_double[4][15] , \tmp_A_neg_double[4][14] , 
        \tmp_A_neg_double[4][13] , \tmp_A_neg_double[4][12] , 
        \tmp_A_neg_double[4][11] , \tmp_A_neg_double[4][10] , A[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(B[9:7]), .Y({
        \out_mux[4][31] , \out_mux[4][30] , \out_mux[4][29] , \out_mux[4][28] , 
        \out_mux[4][27] , \out_mux[4][26] , \out_mux[4][25] , \out_mux[4][24] , 
        \out_mux[4][23] , \out_mux[4][22] , \out_mux[4][21] , \out_mux[4][20] , 
        \out_mux[4][19] , \out_mux[4][18] , \out_mux[4][17] , \out_mux[4][16] , 
        \out_mux[4][15] , \out_mux[4][14] , \out_mux[4][13] , \out_mux[4][12] , 
        \out_mux[4][11] , \out_mux[4][10] , \out_mux[4][9] , \out_mux[4][8] , 
        \out_mux[4][7] , \out_mux[4][6] , \out_mux[4][5] , \out_mux[4][4] , 
        \out_mux[4][3] , \out_mux[4][2] , \out_mux[4][1] , \out_mux[4][0] })
         );
  P4adder_N32_PowerN5_4 sum_4 ( .A({\out_mux[4][31] , \out_mux[4][30] , 
        \out_mux[4][29] , \out_mux[4][28] , \out_mux[4][27] , \out_mux[4][26] , 
        \out_mux[4][25] , \out_mux[4][24] , \out_mux[4][23] , \out_mux[4][22] , 
        \out_mux[4][21] , \out_mux[4][20] , \out_mux[4][19] , \out_mux[4][18] , 
        \out_mux[4][17] , \out_mux[4][16] , \out_mux[4][15] , \out_mux[4][14] , 
        \out_mux[4][13] , \out_mux[4][12] , \out_mux[4][11] , \out_mux[4][10] , 
        \out_mux[4][9] , \out_mux[4][8] , \out_mux[4][7] , \out_mux[4][6] , 
        \out_mux[4][5] , \out_mux[4][4] , \out_mux[4][3] , \out_mux[4][2] , 
        \out_mux[4][1] , \out_mux[4][0] }), .B({\out_sum[2][31] , 
        \out_sum[2][30] , \out_sum[2][29] , \out_sum[2][28] , \out_sum[2][27] , 
        \out_sum[2][26] , \out_sum[2][25] , \out_sum[2][24] , \out_sum[2][23] , 
        \out_sum[2][22] , \out_sum[2][21] , \out_sum[2][20] , \out_sum[2][19] , 
        \out_sum[2][18] , \out_sum[2][17] , \out_sum[2][16] , \out_sum[2][15] , 
        \out_sum[2][14] , \out_sum[2][13] , \out_sum[2][12] , \out_sum[2][11] , 
        \out_sum[2][10] , \out_sum[2][9] , \out_sum[2][8] , \out_sum[2][7] , 
        \out_sum[2][6] , \out_sum[2][5] , \out_sum[2][4] , \out_sum[2][3] , 
        \out_sum[2][2] , \out_sum[2][1] , \out_sum[2][0] }), .Ci(1'b0), .S({
        \out_sum[3][31] , \out_sum[3][30] , \out_sum[3][29] , \out_sum[3][28] , 
        \out_sum[3][27] , \out_sum[3][26] , \out_sum[3][25] , \out_sum[3][24] , 
        \out_sum[3][23] , \out_sum[3][22] , \out_sum[3][21] , \out_sum[3][20] , 
        \out_sum[3][19] , \out_sum[3][18] , \out_sum[3][17] , \out_sum[3][16] , 
        \out_sum[3][15] , \out_sum[3][14] , \out_sum[3][13] , \out_sum[3][12] , 
        \out_sum[3][11] , \out_sum[3][10] , \out_sum[3][9] , \out_sum[3][8] , 
        \out_sum[3][7] , \out_sum[3][6] , \out_sum[3][5] , \out_sum[3][4] , 
        \out_sum[3][3] , \out_sum[3][2] , \out_sum[3][1] , \out_sum[3][0] })
         );
  booth_mux_generic_N32_3 Muxes_5 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n66, n65, n65, n65, n65, n65, n65, A[14:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[5][31] , \tmp_A_neg[5][30] , \tmp_A_neg[5][29] , 
        \tmp_A_neg[5][28] , \tmp_A_neg[5][27] , \tmp_A_neg[5][26] , 
        \tmp_A_neg[5][25] , \tmp_A_neg[5][24] , \tmp_A_neg[5][23] , 
        \tmp_A_neg[5][22] , \tmp_A_neg[5][21] , \tmp_A_neg[5][20] , 
        \tmp_A_neg[5][19] , \tmp_A_neg[5][18] , \tmp_A_neg[5][17] , 
        \tmp_A_neg[5][16] , \tmp_A_neg[5][15] , \tmp_A_neg[5][14] , 
        \tmp_A_neg[5][13] , \tmp_A_neg[5][12] , \tmp_A_neg[5][11] , 
        \tmp_A_neg[5][10] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A_double({n65, n65, n65, n65, n65, n65, A[14:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .A_neg_double({\tmp_A_neg_double[5][31] , \tmp_A_neg_double[5][30] , 
        \tmp_A_neg_double[5][29] , \tmp_A_neg_double[5][28] , 
        \tmp_A_neg_double[5][27] , \tmp_A_neg_double[5][26] , 
        \tmp_A_neg_double[5][25] , \tmp_A_neg_double[5][24] , 
        \tmp_A_neg_double[5][23] , \tmp_A_neg_double[5][22] , 
        \tmp_A_neg_double[5][21] , \tmp_A_neg_double[5][20] , 
        \tmp_A_neg_double[5][19] , \tmp_A_neg_double[5][18] , 
        \tmp_A_neg_double[5][17] , \tmp_A_neg_double[5][16] , 
        \tmp_A_neg_double[5][15] , \tmp_A_neg_double[5][14] , 
        \tmp_A_neg_double[5][13] , \tmp_A_neg_double[5][12] , 
        \tmp_A_neg_double[5][11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .SEL(B[11:9]), .Y({\out_mux[5][31] , 
        \out_mux[5][30] , \out_mux[5][29] , \out_mux[5][28] , \out_mux[5][27] , 
        \out_mux[5][26] , \out_mux[5][25] , \out_mux[5][24] , \out_mux[5][23] , 
        \out_mux[5][22] , \out_mux[5][21] , \out_mux[5][20] , \out_mux[5][19] , 
        \out_mux[5][18] , \out_mux[5][17] , \out_mux[5][16] , \out_mux[5][15] , 
        \out_mux[5][14] , \out_mux[5][13] , \out_mux[5][12] , \out_mux[5][11] , 
        \out_mux[5][10] , \out_mux[5][9] , \out_mux[5][8] , \out_mux[5][7] , 
        \out_mux[5][6] , \out_mux[5][5] , \out_mux[5][4] , \out_mux[5][3] , 
        \out_mux[5][2] , \out_mux[5][1] , \out_mux[5][0] }) );
  P4adder_N32_PowerN5_3 sum_5 ( .A({\out_mux[5][31] , \out_mux[5][30] , 
        \out_mux[5][29] , \out_mux[5][28] , \out_mux[5][27] , \out_mux[5][26] , 
        \out_mux[5][25] , \out_mux[5][24] , \out_mux[5][23] , \out_mux[5][22] , 
        \out_mux[5][21] , \out_mux[5][20] , \out_mux[5][19] , \out_mux[5][18] , 
        \out_mux[5][17] , \out_mux[5][16] , \out_mux[5][15] , \out_mux[5][14] , 
        \out_mux[5][13] , \out_mux[5][12] , \out_mux[5][11] , \out_mux[5][10] , 
        \out_mux[5][9] , \out_mux[5][8] , \out_mux[5][7] , \out_mux[5][6] , 
        \out_mux[5][5] , \out_mux[5][4] , \out_mux[5][3] , \out_mux[5][2] , 
        \out_mux[5][1] , \out_mux[5][0] }), .B({\out_sum[3][31] , 
        \out_sum[3][30] , \out_sum[3][29] , \out_sum[3][28] , \out_sum[3][27] , 
        \out_sum[3][26] , \out_sum[3][25] , \out_sum[3][24] , \out_sum[3][23] , 
        \out_sum[3][22] , \out_sum[3][21] , \out_sum[3][20] , \out_sum[3][19] , 
        \out_sum[3][18] , \out_sum[3][17] , \out_sum[3][16] , \out_sum[3][15] , 
        \out_sum[3][14] , \out_sum[3][13] , \out_sum[3][12] , \out_sum[3][11] , 
        \out_sum[3][10] , \out_sum[3][9] , \out_sum[3][8] , \out_sum[3][7] , 
        \out_sum[3][6] , \out_sum[3][5] , \out_sum[3][4] , \out_sum[3][3] , 
        \out_sum[3][2] , \out_sum[3][1] , \out_sum[3][0] }), .Ci(1'b0), .S({
        \out_sum[4][31] , \out_sum[4][30] , \out_sum[4][29] , \out_sum[4][28] , 
        \out_sum[4][27] , \out_sum[4][26] , \out_sum[4][25] , \out_sum[4][24] , 
        \out_sum[4][23] , \out_sum[4][22] , \out_sum[4][21] , \out_sum[4][20] , 
        \out_sum[4][19] , \out_sum[4][18] , \out_sum[4][17] , \out_sum[4][16] , 
        \out_sum[4][15] , \out_sum[4][14] , \out_sum[4][13] , \out_sum[4][12] , 
        \out_sum[4][11] , \out_sum[4][10] , \out_sum[4][9] , \out_sum[4][8] , 
        \out_sum[4][7] , \out_sum[4][6] , \out_sum[4][5] , \out_sum[4][4] , 
        \out_sum[4][3] , \out_sum[4][2] , \out_sum[4][1] , \out_sum[4][0] })
         );
  booth_mux_generic_N32_2 Muxes_6 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n66, n66, n66, n66, n66, A[14:0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[6][31] , \tmp_A_neg[6][30] , \tmp_A_neg[6][29] , 
        \tmp_A_neg[6][28] , \tmp_A_neg[6][27] , \tmp_A_neg[6][26] , 
        \tmp_A_neg[6][25] , \tmp_A_neg[6][24] , \tmp_A_neg[6][23] , 
        \tmp_A_neg[6][22] , \tmp_A_neg[6][21] , \tmp_A_neg[6][20] , 
        \tmp_A_neg[6][19] , \tmp_A_neg[6][18] , \tmp_A_neg[6][17] , 
        \tmp_A_neg[6][16] , \tmp_A_neg[6][15] , \tmp_A_neg[6][14] , 
        \tmp_A_neg[6][13] , A[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_double({n66, n66, n66, n66, A[14:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .A_neg_double({\tmp_A_neg_double[6][31] , 
        \tmp_A_neg_double[6][30] , \tmp_A_neg_double[6][29] , 
        \tmp_A_neg_double[6][28] , \tmp_A_neg_double[6][27] , 
        \tmp_A_neg_double[6][26] , \tmp_A_neg_double[6][25] , 
        \tmp_A_neg_double[6][24] , \tmp_A_neg_double[6][23] , 
        \tmp_A_neg_double[6][22] , \tmp_A_neg_double[6][21] , 
        \tmp_A_neg_double[6][20] , \tmp_A_neg_double[6][19] , 
        \tmp_A_neg_double[6][18] , \tmp_A_neg_double[6][17] , 
        \tmp_A_neg_double[6][16] , \tmp_A_neg_double[6][15] , 
        \tmp_A_neg_double[6][14] , A[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(B[13:11]), .Y({
        \out_mux[6][31] , \out_mux[6][30] , \out_mux[6][29] , \out_mux[6][28] , 
        \out_mux[6][27] , \out_mux[6][26] , \out_mux[6][25] , \out_mux[6][24] , 
        \out_mux[6][23] , \out_mux[6][22] , \out_mux[6][21] , \out_mux[6][20] , 
        \out_mux[6][19] , \out_mux[6][18] , \out_mux[6][17] , \out_mux[6][16] , 
        \out_mux[6][15] , \out_mux[6][14] , \out_mux[6][13] , \out_mux[6][12] , 
        \out_mux[6][11] , \out_mux[6][10] , \out_mux[6][9] , \out_mux[6][8] , 
        \out_mux[6][7] , \out_mux[6][6] , \out_mux[6][5] , \out_mux[6][4] , 
        \out_mux[6][3] , \out_mux[6][2] , \out_mux[6][1] , \out_mux[6][0] })
         );
  P4adder_N32_PowerN5_2 sum_6 ( .A({\out_mux[6][31] , \out_mux[6][30] , 
        \out_mux[6][29] , \out_mux[6][28] , \out_mux[6][27] , \out_mux[6][26] , 
        \out_mux[6][25] , \out_mux[6][24] , \out_mux[6][23] , \out_mux[6][22] , 
        \out_mux[6][21] , \out_mux[6][20] , \out_mux[6][19] , \out_mux[6][18] , 
        \out_mux[6][17] , \out_mux[6][16] , \out_mux[6][15] , \out_mux[6][14] , 
        \out_mux[6][13] , \out_mux[6][12] , \out_mux[6][11] , \out_mux[6][10] , 
        \out_mux[6][9] , \out_mux[6][8] , \out_mux[6][7] , \out_mux[6][6] , 
        \out_mux[6][5] , \out_mux[6][4] , \out_mux[6][3] , \out_mux[6][2] , 
        \out_mux[6][1] , \out_mux[6][0] }), .B({\out_sum[4][31] , 
        \out_sum[4][30] , \out_sum[4][29] , \out_sum[4][28] , \out_sum[4][27] , 
        \out_sum[4][26] , \out_sum[4][25] , \out_sum[4][24] , \out_sum[4][23] , 
        \out_sum[4][22] , \out_sum[4][21] , \out_sum[4][20] , \out_sum[4][19] , 
        \out_sum[4][18] , \out_sum[4][17] , \out_sum[4][16] , \out_sum[4][15] , 
        \out_sum[4][14] , \out_sum[4][13] , \out_sum[4][12] , \out_sum[4][11] , 
        \out_sum[4][10] , \out_sum[4][9] , \out_sum[4][8] , \out_sum[4][7] , 
        \out_sum[4][6] , \out_sum[4][5] , \out_sum[4][4] , \out_sum[4][3] , 
        \out_sum[4][2] , \out_sum[4][1] , \out_sum[4][0] }), .Ci(1'b0), .S({
        \out_sum[5][31] , \out_sum[5][30] , \out_sum[5][29] , \out_sum[5][28] , 
        \out_sum[5][27] , \out_sum[5][26] , \out_sum[5][25] , \out_sum[5][24] , 
        \out_sum[5][23] , \out_sum[5][22] , \out_sum[5][21] , \out_sum[5][20] , 
        \out_sum[5][19] , \out_sum[5][18] , \out_sum[5][17] , \out_sum[5][16] , 
        \out_sum[5][15] , \out_sum[5][14] , \out_sum[5][13] , \out_sum[5][12] , 
        \out_sum[5][11] , \out_sum[5][10] , \out_sum[5][9] , \out_sum[5][8] , 
        \out_sum[5][7] , \out_sum[5][6] , \out_sum[5][5] , \out_sum[5][4] , 
        \out_sum[5][3] , \out_sum[5][2] , \out_sum[5][1] , \out_sum[5][0] })
         );
  booth_mux_generic_N32_1 Muxes_7 ( .Zero({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .A({n67, n67, n66, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg({
        \tmp_A_neg[7][31] , \tmp_A_neg[7][30] , \tmp_A_neg[7][29] , 
        \tmp_A_neg[7][28] , \tmp_A_neg[7][27] , \tmp_A_neg[7][26] , 
        \tmp_A_neg[7][25] , \tmp_A_neg[7][24] , \tmp_A_neg[7][23] , 
        \tmp_A_neg[7][22] , \tmp_A_neg[7][21] , \tmp_A_neg[7][20] , 
        \tmp_A_neg[7][19] , \tmp_A_neg[7][18] , \tmp_A_neg[7][17] , 
        \tmp_A_neg[7][16] , \tmp_A_neg[7][15] , A[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .A_double({n66, n66, A[14:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_neg_double({
        \tmp_A_neg_double[7][31] , \tmp_A_neg_double[7][30] , 
        \tmp_A_neg_double[7][29] , \tmp_A_neg_double[7][28] , 
        \tmp_A_neg_double[7][27] , \tmp_A_neg_double[7][26] , 
        \tmp_A_neg_double[7][25] , \tmp_A_neg_double[7][24] , 
        \tmp_A_neg_double[7][23] , \tmp_A_neg_double[7][22] , 
        \tmp_A_neg_double[7][21] , \tmp_A_neg_double[7][20] , 
        \tmp_A_neg_double[7][19] , \tmp_A_neg_double[7][18] , 
        \tmp_A_neg_double[7][17] , \tmp_A_neg_double[7][16] , A[0], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SEL(B[15:13]), .Y({\out_mux[7][31] , \out_mux[7][30] , 
        \out_mux[7][29] , \out_mux[7][28] , \out_mux[7][27] , \out_mux[7][26] , 
        \out_mux[7][25] , \out_mux[7][24] , \out_mux[7][23] , \out_mux[7][22] , 
        \out_mux[7][21] , \out_mux[7][20] , \out_mux[7][19] , \out_mux[7][18] , 
        \out_mux[7][17] , \out_mux[7][16] , \out_mux[7][15] , \out_mux[7][14] , 
        \out_mux[7][13] , \out_mux[7][12] , \out_mux[7][11] , \out_mux[7][10] , 
        \out_mux[7][9] , \out_mux[7][8] , \out_mux[7][7] , \out_mux[7][6] , 
        \out_mux[7][5] , \out_mux[7][4] , \out_mux[7][3] , \out_mux[7][2] , 
        \out_mux[7][1] , \out_mux[7][0] }) );
  P4adder_N32_PowerN5_1 sum_7 ( .A({\out_mux[7][31] , \out_mux[7][30] , 
        \out_mux[7][29] , \out_mux[7][28] , \out_mux[7][27] , \out_mux[7][26] , 
        \out_mux[7][25] , \out_mux[7][24] , \out_mux[7][23] , \out_mux[7][22] , 
        \out_mux[7][21] , \out_mux[7][20] , \out_mux[7][19] , \out_mux[7][18] , 
        \out_mux[7][17] , \out_mux[7][16] , \out_mux[7][15] , \out_mux[7][14] , 
        \out_mux[7][13] , \out_mux[7][12] , \out_mux[7][11] , \out_mux[7][10] , 
        \out_mux[7][9] , \out_mux[7][8] , \out_mux[7][7] , \out_mux[7][6] , 
        \out_mux[7][5] , \out_mux[7][4] , \out_mux[7][3] , \out_mux[7][2] , 
        \out_mux[7][1] , \out_mux[7][0] }), .B({\out_sum[5][31] , 
        \out_sum[5][30] , \out_sum[5][29] , \out_sum[5][28] , \out_sum[5][27] , 
        \out_sum[5][26] , \out_sum[5][25] , \out_sum[5][24] , \out_sum[5][23] , 
        \out_sum[5][22] , \out_sum[5][21] , \out_sum[5][20] , \out_sum[5][19] , 
        \out_sum[5][18] , \out_sum[5][17] , \out_sum[5][16] , \out_sum[5][15] , 
        \out_sum[5][14] , \out_sum[5][13] , \out_sum[5][12] , \out_sum[5][11] , 
        \out_sum[5][10] , \out_sum[5][9] , \out_sum[5][8] , \out_sum[5][7] , 
        \out_sum[5][6] , \out_sum[5][5] , \out_sum[5][4] , \out_sum[5][3] , 
        \out_sum[5][2] , \out_sum[5][1] , \out_sum[5][0] }), .Ci(1'b0), .S(Res) );
  boothmul_Nbit16_DW01_inc_4 add_83_2_C132_G6 ( .A({n77, n76, n76, n74, n72, 
        n72, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, n41, n56, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .SUM({\tmp_A_neg_double[5][31] , \tmp_A_neg_double[5][30] , 
        \tmp_A_neg_double[5][29] , \tmp_A_neg_double[5][28] , 
        \tmp_A_neg_double[5][27] , \tmp_A_neg_double[5][26] , 
        \tmp_A_neg_double[5][25] , \tmp_A_neg_double[5][24] , 
        \tmp_A_neg_double[5][23] , \tmp_A_neg_double[5][22] , 
        \tmp_A_neg_double[5][21] , \tmp_A_neg_double[5][20] , 
        \tmp_A_neg_double[5][19] , \tmp_A_neg_double[5][18] , 
        \tmp_A_neg_double[5][17] , \tmp_A_neg_double[5][16] , 
        \tmp_A_neg_double[5][15] , \tmp_A_neg_double[5][14] , 
        \tmp_A_neg_double[5][13] , \tmp_A_neg_double[5][12] , 
        \tmp_A_neg_double[5][11] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10}) );
  boothmul_Nbit16_DW01_inc_5 add_83_2_C130_G6 ( .A({n74, n76, n73, n71, n73, 
        n72, n71, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, n41, 
        n56, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .SUM({\tmp_A_neg[5][31] , \tmp_A_neg[5][30] , \tmp_A_neg[5][29] , 
        \tmp_A_neg[5][28] , \tmp_A_neg[5][27] , \tmp_A_neg[5][26] , 
        \tmp_A_neg[5][25] , \tmp_A_neg[5][24] , \tmp_A_neg[5][23] , 
        \tmp_A_neg[5][22] , \tmp_A_neg[5][21] , \tmp_A_neg[5][20] , 
        \tmp_A_neg[5][19] , \tmp_A_neg[5][18] , \tmp_A_neg[5][17] , 
        \tmp_A_neg[5][16] , \tmp_A_neg[5][15] , \tmp_A_neg[5][14] , 
        \tmp_A_neg[5][13] , \tmp_A_neg[5][12] , \tmp_A_neg[5][11] , 
        \tmp_A_neg[5][10] , SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20}) );
  HA_X1 \add_83_2_C132_G8/U1_1_16  ( .A(n41), .B(n56), .CO(
        \add_83_2_C132_G8/carry[17] ), .S(\tmp_A_neg_double[7][16] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_17  ( .A(N13), .B(\add_83_2_C132_G8/carry[17] ), 
        .CO(\add_83_2_C132_G8/carry[18] ), .S(\tmp_A_neg_double[7][17] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_18  ( .A(N12), .B(\add_83_2_C132_G8/carry[18] ), 
        .CO(\add_83_2_C132_G8/carry[19] ), .S(\tmp_A_neg_double[7][18] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_19  ( .A(N11), .B(\add_83_2_C132_G8/carry[19] ), 
        .CO(\add_83_2_C132_G8/carry[20] ), .S(\tmp_A_neg_double[7][19] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_20  ( .A(N10), .B(\add_83_2_C132_G8/carry[20] ), 
        .CO(\add_83_2_C132_G8/carry[21] ), .S(\tmp_A_neg_double[7][20] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_21  ( .A(N9), .B(\add_83_2_C132_G8/carry[21] ), 
        .CO(\add_83_2_C132_G8/carry[22] ), .S(\tmp_A_neg_double[7][21] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_22  ( .A(N8), .B(\add_83_2_C132_G8/carry[22] ), 
        .CO(\add_83_2_C132_G8/carry[23] ), .S(\tmp_A_neg_double[7][22] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_23  ( .A(N7), .B(\add_83_2_C132_G8/carry[23] ), 
        .CO(\add_83_2_C132_G8/carry[24] ), .S(\tmp_A_neg_double[7][23] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_24  ( .A(N6), .B(\add_83_2_C132_G8/carry[24] ), 
        .CO(\add_83_2_C132_G8/carry[25] ), .S(\tmp_A_neg_double[7][24] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_25  ( .A(N5), .B(\add_83_2_C132_G8/carry[25] ), 
        .CO(\add_83_2_C132_G8/carry[26] ), .S(\tmp_A_neg_double[7][25] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_26  ( .A(N4), .B(\add_83_2_C132_G8/carry[26] ), 
        .CO(\add_83_2_C132_G8/carry[27] ), .S(\tmp_A_neg_double[7][26] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_27  ( .A(N3), .B(\add_83_2_C132_G8/carry[27] ), 
        .CO(\add_83_2_C132_G8/carry[28] ), .S(\tmp_A_neg_double[7][27] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_28  ( .A(N2), .B(\add_83_2_C132_G8/carry[28] ), 
        .CO(\add_83_2_C132_G8/carry[29] ), .S(\tmp_A_neg_double[7][28] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_29  ( .A(N1), .B(\add_83_2_C132_G8/carry[29] ), 
        .CO(\add_83_2_C132_G8/carry[30] ), .S(\tmp_A_neg_double[7][29] ) );
  HA_X1 \add_83_2_C132_G8/U1_1_30  ( .A(n75), .B(\add_83_2_C132_G8/carry[30] ), 
        .CO(\add_83_2_C132_G8/carry[31] ), .S(\tmp_A_neg_double[7][30] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_15  ( .A(n41), .B(n56), .CO(
        \add_83_2_C130_G8/carry[16] ), .S(\tmp_A_neg[7][15] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_16  ( .A(N13), .B(\add_83_2_C130_G8/carry[16] ), 
        .CO(\add_83_2_C130_G8/carry[17] ), .S(\tmp_A_neg[7][16] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_17  ( .A(N12), .B(\add_83_2_C130_G8/carry[17] ), 
        .CO(\add_83_2_C130_G8/carry[18] ), .S(\tmp_A_neg[7][17] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_18  ( .A(N11), .B(\add_83_2_C130_G8/carry[18] ), 
        .CO(\add_83_2_C130_G8/carry[19] ), .S(\tmp_A_neg[7][18] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_19  ( .A(N10), .B(\add_83_2_C130_G8/carry[19] ), 
        .CO(\add_83_2_C130_G8/carry[20] ), .S(\tmp_A_neg[7][19] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_20  ( .A(N9), .B(\add_83_2_C130_G8/carry[20] ), 
        .CO(\add_83_2_C130_G8/carry[21] ), .S(\tmp_A_neg[7][20] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_21  ( .A(N8), .B(\add_83_2_C130_G8/carry[21] ), 
        .CO(\add_83_2_C130_G8/carry[22] ), .S(\tmp_A_neg[7][21] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_22  ( .A(N7), .B(\add_83_2_C130_G8/carry[22] ), 
        .CO(\add_83_2_C130_G8/carry[23] ), .S(\tmp_A_neg[7][22] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_23  ( .A(N6), .B(\add_83_2_C130_G8/carry[23] ), 
        .CO(\add_83_2_C130_G8/carry[24] ), .S(\tmp_A_neg[7][23] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_24  ( .A(N5), .B(\add_83_2_C130_G8/carry[24] ), 
        .CO(\add_83_2_C130_G8/carry[25] ), .S(\tmp_A_neg[7][24] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_25  ( .A(N4), .B(\add_83_2_C130_G8/carry[25] ), 
        .CO(\add_83_2_C130_G8/carry[26] ), .S(\tmp_A_neg[7][25] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_26  ( .A(N3), .B(\add_83_2_C130_G8/carry[26] ), 
        .CO(\add_83_2_C130_G8/carry[27] ), .S(\tmp_A_neg[7][26] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_27  ( .A(N2), .B(\add_83_2_C130_G8/carry[27] ), 
        .CO(\add_83_2_C130_G8/carry[28] ), .S(\tmp_A_neg[7][27] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_28  ( .A(N1), .B(\add_83_2_C130_G8/carry[28] ), 
        .CO(\add_83_2_C130_G8/carry[29] ), .S(\tmp_A_neg[7][28] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_29  ( .A(n75), .B(\add_83_2_C130_G8/carry[29] ), 
        .CO(\add_83_2_C130_G8/carry[30] ), .S(\tmp_A_neg[7][29] ) );
  HA_X1 \add_83_2_C130_G8/U1_1_30  ( .A(n75), .B(\add_83_2_C130_G8/carry[30] ), 
        .CO(\add_83_2_C130_G8/carry[31] ), .S(\tmp_A_neg[7][30] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_14  ( .A(n41), .B(n56), .CO(
        \add_83_2_C132_G7/carry[15] ), .S(\tmp_A_neg_double[6][14] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_15  ( .A(N13), .B(\add_83_2_C132_G7/carry[15] ), 
        .CO(\add_83_2_C132_G7/carry[16] ), .S(\tmp_A_neg_double[6][15] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_16  ( .A(N12), .B(\add_83_2_C132_G7/carry[16] ), 
        .CO(\add_83_2_C132_G7/carry[17] ), .S(\tmp_A_neg_double[6][16] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_17  ( .A(N11), .B(\add_83_2_C132_G7/carry[17] ), 
        .CO(\add_83_2_C132_G7/carry[18] ), .S(\tmp_A_neg_double[6][17] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_18  ( .A(N10), .B(\add_83_2_C132_G7/carry[18] ), 
        .CO(\add_83_2_C132_G7/carry[19] ), .S(\tmp_A_neg_double[6][18] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_19  ( .A(N9), .B(\add_83_2_C132_G7/carry[19] ), 
        .CO(\add_83_2_C132_G7/carry[20] ), .S(\tmp_A_neg_double[6][19] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_20  ( .A(N8), .B(\add_83_2_C132_G7/carry[20] ), 
        .CO(\add_83_2_C132_G7/carry[21] ), .S(\tmp_A_neg_double[6][20] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_21  ( .A(N7), .B(\add_83_2_C132_G7/carry[21] ), 
        .CO(\add_83_2_C132_G7/carry[22] ), .S(\tmp_A_neg_double[6][21] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_22  ( .A(N6), .B(\add_83_2_C132_G7/carry[22] ), 
        .CO(\add_83_2_C132_G7/carry[23] ), .S(\tmp_A_neg_double[6][22] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_23  ( .A(N5), .B(\add_83_2_C132_G7/carry[23] ), 
        .CO(\add_83_2_C132_G7/carry[24] ), .S(\tmp_A_neg_double[6][23] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_24  ( .A(N4), .B(\add_83_2_C132_G7/carry[24] ), 
        .CO(\add_83_2_C132_G7/carry[25] ), .S(\tmp_A_neg_double[6][24] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_25  ( .A(N3), .B(\add_83_2_C132_G7/carry[25] ), 
        .CO(\add_83_2_C132_G7/carry[26] ), .S(\tmp_A_neg_double[6][25] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_26  ( .A(N2), .B(\add_83_2_C132_G7/carry[26] ), 
        .CO(\add_83_2_C132_G7/carry[27] ), .S(\tmp_A_neg_double[6][26] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_27  ( .A(N1), .B(\add_83_2_C132_G7/carry[27] ), 
        .CO(\add_83_2_C132_G7/carry[28] ), .S(\tmp_A_neg_double[6][27] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_28  ( .A(n75), .B(\add_83_2_C132_G7/carry[28] ), 
        .CO(\add_83_2_C132_G7/carry[29] ), .S(\tmp_A_neg_double[6][28] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_29  ( .A(n76), .B(\add_83_2_C132_G7/carry[29] ), 
        .CO(\add_83_2_C132_G7/carry[30] ), .S(\tmp_A_neg_double[6][29] ) );
  HA_X1 \add_83_2_C132_G7/U1_1_30  ( .A(n75), .B(\add_83_2_C132_G7/carry[30] ), 
        .CO(\add_83_2_C132_G7/carry[31] ), .S(\tmp_A_neg_double[6][30] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_13  ( .A(n41), .B(n56), .CO(
        \add_83_2_C130_G7/carry[14] ), .S(\tmp_A_neg[6][13] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_14  ( .A(N13), .B(\add_83_2_C130_G7/carry[14] ), 
        .CO(\add_83_2_C130_G7/carry[15] ), .S(\tmp_A_neg[6][14] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_15  ( .A(N12), .B(\add_83_2_C130_G7/carry[15] ), 
        .CO(\add_83_2_C130_G7/carry[16] ), .S(\tmp_A_neg[6][15] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_16  ( .A(N11), .B(\add_83_2_C130_G7/carry[16] ), 
        .CO(\add_83_2_C130_G7/carry[17] ), .S(\tmp_A_neg[6][16] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_17  ( .A(N10), .B(\add_83_2_C130_G7/carry[17] ), 
        .CO(\add_83_2_C130_G7/carry[18] ), .S(\tmp_A_neg[6][17] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_18  ( .A(N9), .B(\add_83_2_C130_G7/carry[18] ), 
        .CO(\add_83_2_C130_G7/carry[19] ), .S(\tmp_A_neg[6][18] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_19  ( .A(N8), .B(\add_83_2_C130_G7/carry[19] ), 
        .CO(\add_83_2_C130_G7/carry[20] ), .S(\tmp_A_neg[6][19] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_20  ( .A(N7), .B(\add_83_2_C130_G7/carry[20] ), 
        .CO(\add_83_2_C130_G7/carry[21] ), .S(\tmp_A_neg[6][20] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_21  ( .A(N6), .B(\add_83_2_C130_G7/carry[21] ), 
        .CO(\add_83_2_C130_G7/carry[22] ), .S(\tmp_A_neg[6][21] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_22  ( .A(N5), .B(\add_83_2_C130_G7/carry[22] ), 
        .CO(\add_83_2_C130_G7/carry[23] ), .S(\tmp_A_neg[6][22] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_23  ( .A(N4), .B(\add_83_2_C130_G7/carry[23] ), 
        .CO(\add_83_2_C130_G7/carry[24] ), .S(\tmp_A_neg[6][23] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_24  ( .A(N3), .B(\add_83_2_C130_G7/carry[24] ), 
        .CO(\add_83_2_C130_G7/carry[25] ), .S(\tmp_A_neg[6][24] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_25  ( .A(N2), .B(\add_83_2_C130_G7/carry[25] ), 
        .CO(\add_83_2_C130_G7/carry[26] ), .S(\tmp_A_neg[6][25] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_26  ( .A(N1), .B(\add_83_2_C130_G7/carry[26] ), 
        .CO(\add_83_2_C130_G7/carry[27] ), .S(\tmp_A_neg[6][26] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_27  ( .A(n74), .B(\add_83_2_C130_G7/carry[27] ), 
        .CO(\add_83_2_C130_G7/carry[28] ), .S(\tmp_A_neg[6][27] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_28  ( .A(n74), .B(\add_83_2_C130_G7/carry[28] ), 
        .CO(\add_83_2_C130_G7/carry[29] ), .S(\tmp_A_neg[6][28] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_29  ( .A(n76), .B(\add_83_2_C130_G7/carry[29] ), 
        .CO(\add_83_2_C130_G7/carry[30] ), .S(\tmp_A_neg[6][29] ) );
  HA_X1 \add_83_2_C130_G7/U1_1_30  ( .A(n74), .B(\add_83_2_C130_G7/carry[30] ), 
        .CO(\add_83_2_C130_G7/carry[31] ), .S(\tmp_A_neg[6][30] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_10  ( .A(n41), .B(n56), .CO(
        \add_83_2_C132_G5/carry[11] ), .S(\tmp_A_neg_double[4][10] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_11  ( .A(N13), .B(\add_83_2_C132_G5/carry[11] ), 
        .CO(\add_83_2_C132_G5/carry[12] ), .S(\tmp_A_neg_double[4][11] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_12  ( .A(N12), .B(\add_83_2_C132_G5/carry[12] ), 
        .CO(\add_83_2_C132_G5/carry[13] ), .S(\tmp_A_neg_double[4][12] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_13  ( .A(N11), .B(\add_83_2_C132_G5/carry[13] ), 
        .CO(\add_83_2_C132_G5/carry[14] ), .S(\tmp_A_neg_double[4][13] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_14  ( .A(N10), .B(\add_83_2_C132_G5/carry[14] ), 
        .CO(\add_83_2_C132_G5/carry[15] ), .S(\tmp_A_neg_double[4][14] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_15  ( .A(N9), .B(\add_83_2_C132_G5/carry[15] ), 
        .CO(\add_83_2_C132_G5/carry[16] ), .S(\tmp_A_neg_double[4][15] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_16  ( .A(N8), .B(\add_83_2_C132_G5/carry[16] ), 
        .CO(\add_83_2_C132_G5/carry[17] ), .S(\tmp_A_neg_double[4][16] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_17  ( .A(N7), .B(\add_83_2_C132_G5/carry[17] ), 
        .CO(\add_83_2_C132_G5/carry[18] ), .S(\tmp_A_neg_double[4][17] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_18  ( .A(N6), .B(\add_83_2_C132_G5/carry[18] ), 
        .CO(\add_83_2_C132_G5/carry[19] ), .S(\tmp_A_neg_double[4][18] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_19  ( .A(N5), .B(\add_83_2_C132_G5/carry[19] ), 
        .CO(\add_83_2_C132_G5/carry[20] ), .S(\tmp_A_neg_double[4][19] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_20  ( .A(N4), .B(\add_83_2_C132_G5/carry[20] ), 
        .CO(\add_83_2_C132_G5/carry[21] ), .S(\tmp_A_neg_double[4][20] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_21  ( .A(N3), .B(\add_83_2_C132_G5/carry[21] ), 
        .CO(\add_83_2_C132_G5/carry[22] ), .S(\tmp_A_neg_double[4][21] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_22  ( .A(N2), .B(\add_83_2_C132_G5/carry[22] ), 
        .CO(\add_83_2_C132_G5/carry[23] ), .S(\tmp_A_neg_double[4][22] ) );
  HA_X1 \add_83_2_C132_G5/U1_1_23  ( .A(N1), .B(\add_83_2_C132_G5/carry[23] ), 
        .CO(\add_83_2_C132_G5/carry[24] ), .S(\tmp_A_neg_double[4][23] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_9  ( .A(n41), .B(n56), .CO(
        \add_83_2_C130_G5/carry[10] ), .S(\tmp_A_neg[4][9] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_10  ( .A(N13), .B(\add_83_2_C130_G5/carry[10] ), 
        .CO(\add_83_2_C130_G5/carry[11] ), .S(\tmp_A_neg[4][10] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_11  ( .A(N12), .B(\add_83_2_C130_G5/carry[11] ), 
        .CO(\add_83_2_C130_G5/carry[12] ), .S(\tmp_A_neg[4][11] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_12  ( .A(N11), .B(\add_83_2_C130_G5/carry[12] ), 
        .CO(\add_83_2_C130_G5/carry[13] ), .S(\tmp_A_neg[4][12] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_13  ( .A(N10), .B(\add_83_2_C130_G5/carry[13] ), 
        .CO(\add_83_2_C130_G5/carry[14] ), .S(\tmp_A_neg[4][13] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_14  ( .A(N9), .B(\add_83_2_C130_G5/carry[14] ), 
        .CO(\add_83_2_C130_G5/carry[15] ), .S(\tmp_A_neg[4][14] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_15  ( .A(N8), .B(\add_83_2_C130_G5/carry[15] ), 
        .CO(\add_83_2_C130_G5/carry[16] ), .S(\tmp_A_neg[4][15] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_16  ( .A(N7), .B(\add_83_2_C130_G5/carry[16] ), 
        .CO(\add_83_2_C130_G5/carry[17] ), .S(\tmp_A_neg[4][16] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_17  ( .A(N6), .B(\add_83_2_C130_G5/carry[17] ), 
        .CO(\add_83_2_C130_G5/carry[18] ), .S(\tmp_A_neg[4][17] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_18  ( .A(N5), .B(\add_83_2_C130_G5/carry[18] ), 
        .CO(\add_83_2_C130_G5/carry[19] ), .S(\tmp_A_neg[4][18] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_19  ( .A(N4), .B(\add_83_2_C130_G5/carry[19] ), 
        .CO(\add_83_2_C130_G5/carry[20] ), .S(\tmp_A_neg[4][19] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_20  ( .A(N3), .B(\add_83_2_C130_G5/carry[20] ), 
        .CO(\add_83_2_C130_G5/carry[21] ), .S(\tmp_A_neg[4][20] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_21  ( .A(N2), .B(\add_83_2_C130_G5/carry[21] ), 
        .CO(\add_83_2_C130_G5/carry[22] ), .S(\tmp_A_neg[4][21] ) );
  HA_X1 \add_83_2_C130_G5/U1_1_22  ( .A(N1), .B(\add_83_2_C130_G5/carry[22] ), 
        .CO(\add_83_2_C130_G5/carry[23] ), .S(\tmp_A_neg[4][22] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_8  ( .A(n41), .B(n56), .CO(
        \add_83_2_C132_G4/carry[9] ), .S(\tmp_A_neg_double[3][8] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_9  ( .A(N13), .B(\add_83_2_C132_G4/carry[9] ), 
        .CO(\add_83_2_C132_G4/carry[10] ), .S(\tmp_A_neg_double[3][9] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_10  ( .A(N12), .B(\add_83_2_C132_G4/carry[10] ), 
        .CO(\add_83_2_C132_G4/carry[11] ), .S(\tmp_A_neg_double[3][10] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_11  ( .A(N11), .B(\add_83_2_C132_G4/carry[11] ), 
        .CO(\add_83_2_C132_G4/carry[12] ), .S(\tmp_A_neg_double[3][11] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_12  ( .A(N10), .B(\add_83_2_C132_G4/carry[12] ), 
        .CO(\add_83_2_C132_G4/carry[13] ), .S(\tmp_A_neg_double[3][12] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_13  ( .A(N9), .B(\add_83_2_C132_G4/carry[13] ), 
        .CO(\add_83_2_C132_G4/carry[14] ), .S(\tmp_A_neg_double[3][13] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_14  ( .A(N8), .B(\add_83_2_C132_G4/carry[14] ), 
        .CO(\add_83_2_C132_G4/carry[15] ), .S(\tmp_A_neg_double[3][14] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_15  ( .A(N7), .B(\add_83_2_C132_G4/carry[15] ), 
        .CO(\add_83_2_C132_G4/carry[16] ), .S(\tmp_A_neg_double[3][15] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_16  ( .A(N6), .B(\add_83_2_C132_G4/carry[16] ), 
        .CO(\add_83_2_C132_G4/carry[17] ), .S(\tmp_A_neg_double[3][16] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_17  ( .A(N5), .B(\add_83_2_C132_G4/carry[17] ), 
        .CO(\add_83_2_C132_G4/carry[18] ), .S(\tmp_A_neg_double[3][17] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_18  ( .A(N4), .B(\add_83_2_C132_G4/carry[18] ), 
        .CO(\add_83_2_C132_G4/carry[19] ), .S(\tmp_A_neg_double[3][18] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_19  ( .A(N3), .B(\add_83_2_C132_G4/carry[19] ), 
        .CO(\add_83_2_C132_G4/carry[20] ), .S(\tmp_A_neg_double[3][19] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_20  ( .A(N2), .B(\add_83_2_C132_G4/carry[20] ), 
        .CO(\add_83_2_C132_G4/carry[21] ), .S(\tmp_A_neg_double[3][20] ) );
  HA_X1 \add_83_2_C132_G4/U1_1_21  ( .A(N1), .B(\add_83_2_C132_G4/carry[21] ), 
        .CO(\add_83_2_C132_G4/carry[22] ), .S(\tmp_A_neg_double[3][21] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_7  ( .A(n41), .B(n56), .CO(
        \add_83_2_C130_G4/carry[8] ), .S(\tmp_A_neg[3][7] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_8  ( .A(N13), .B(\add_83_2_C130_G4/carry[8] ), 
        .CO(\add_83_2_C130_G4/carry[9] ), .S(\tmp_A_neg[3][8] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_9  ( .A(N12), .B(\add_83_2_C130_G4/carry[9] ), 
        .CO(\add_83_2_C130_G4/carry[10] ), .S(\tmp_A_neg[3][9] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_10  ( .A(N11), .B(\add_83_2_C130_G4/carry[10] ), 
        .CO(\add_83_2_C130_G4/carry[11] ), .S(\tmp_A_neg[3][10] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_11  ( .A(N10), .B(\add_83_2_C130_G4/carry[11] ), 
        .CO(\add_83_2_C130_G4/carry[12] ), .S(\tmp_A_neg[3][11] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_12  ( .A(N9), .B(\add_83_2_C130_G4/carry[12] ), 
        .CO(\add_83_2_C130_G4/carry[13] ), .S(\tmp_A_neg[3][12] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_13  ( .A(N8), .B(\add_83_2_C130_G4/carry[13] ), 
        .CO(\add_83_2_C130_G4/carry[14] ), .S(\tmp_A_neg[3][13] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_14  ( .A(N7), .B(\add_83_2_C130_G4/carry[14] ), 
        .CO(\add_83_2_C130_G4/carry[15] ), .S(\tmp_A_neg[3][14] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_15  ( .A(N6), .B(\add_83_2_C130_G4/carry[15] ), 
        .CO(\add_83_2_C130_G4/carry[16] ), .S(\tmp_A_neg[3][15] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_16  ( .A(N5), .B(\add_83_2_C130_G4/carry[16] ), 
        .CO(\add_83_2_C130_G4/carry[17] ), .S(\tmp_A_neg[3][16] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_17  ( .A(N4), .B(\add_83_2_C130_G4/carry[17] ), 
        .CO(\add_83_2_C130_G4/carry[18] ), .S(\tmp_A_neg[3][17] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_18  ( .A(N3), .B(\add_83_2_C130_G4/carry[18] ), 
        .CO(\add_83_2_C130_G4/carry[19] ), .S(\tmp_A_neg[3][18] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_19  ( .A(N2), .B(\add_83_2_C130_G4/carry[19] ), 
        .CO(\add_83_2_C130_G4/carry[20] ), .S(\tmp_A_neg[3][19] ) );
  HA_X1 \add_83_2_C130_G4/U1_1_20  ( .A(N1), .B(\add_83_2_C130_G4/carry[20] ), 
        .CO(\add_83_2_C130_G4/carry[21] ), .S(\tmp_A_neg[3][20] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_6  ( .A(n41), .B(n57), .CO(
        \add_83_2_C132_G3/carry[7] ), .S(\tmp_A_neg_double[2][6] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_7  ( .A(N13), .B(\add_83_2_C132_G3/carry[7] ), 
        .CO(\add_83_2_C132_G3/carry[8] ), .S(\tmp_A_neg_double[2][7] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_8  ( .A(N12), .B(\add_83_2_C132_G3/carry[8] ), 
        .CO(\add_83_2_C132_G3/carry[9] ), .S(\tmp_A_neg_double[2][8] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_9  ( .A(N11), .B(\add_83_2_C132_G3/carry[9] ), 
        .CO(\add_83_2_C132_G3/carry[10] ), .S(\tmp_A_neg_double[2][9] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_10  ( .A(N10), .B(\add_83_2_C132_G3/carry[10] ), 
        .CO(\add_83_2_C132_G3/carry[11] ), .S(\tmp_A_neg_double[2][10] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_11  ( .A(N9), .B(\add_83_2_C132_G3/carry[11] ), 
        .CO(\add_83_2_C132_G3/carry[12] ), .S(\tmp_A_neg_double[2][11] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_12  ( .A(N8), .B(\add_83_2_C132_G3/carry[12] ), 
        .CO(\add_83_2_C132_G3/carry[13] ), .S(\tmp_A_neg_double[2][12] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_13  ( .A(N7), .B(\add_83_2_C132_G3/carry[13] ), 
        .CO(\add_83_2_C132_G3/carry[14] ), .S(\tmp_A_neg_double[2][13] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_14  ( .A(N6), .B(\add_83_2_C132_G3/carry[14] ), 
        .CO(\add_83_2_C132_G3/carry[15] ), .S(\tmp_A_neg_double[2][14] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_15  ( .A(N5), .B(\add_83_2_C132_G3/carry[15] ), 
        .CO(\add_83_2_C132_G3/carry[16] ), .S(\tmp_A_neg_double[2][15] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_16  ( .A(N4), .B(\add_83_2_C132_G3/carry[16] ), 
        .CO(\add_83_2_C132_G3/carry[17] ), .S(\tmp_A_neg_double[2][16] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_17  ( .A(N3), .B(\add_83_2_C132_G3/carry[17] ), 
        .CO(\add_83_2_C132_G3/carry[18] ), .S(\tmp_A_neg_double[2][17] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_18  ( .A(N2), .B(\add_83_2_C132_G3/carry[18] ), 
        .CO(\add_83_2_C132_G3/carry[19] ), .S(\tmp_A_neg_double[2][18] ) );
  HA_X1 \add_83_2_C132_G3/U1_1_19  ( .A(N1), .B(\add_83_2_C132_G3/carry[19] ), 
        .CO(\add_83_2_C132_G3/carry[20] ), .S(\tmp_A_neg_double[2][19] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_5  ( .A(n41), .B(n57), .CO(
        \add_83_2_C130_G3/carry[6] ), .S(\tmp_A_neg[2][5] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_6  ( .A(N13), .B(\add_83_2_C130_G3/carry[6] ), 
        .CO(\add_83_2_C130_G3/carry[7] ), .S(\tmp_A_neg[2][6] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_7  ( .A(N12), .B(\add_83_2_C130_G3/carry[7] ), 
        .CO(\add_83_2_C130_G3/carry[8] ), .S(\tmp_A_neg[2][7] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_8  ( .A(N11), .B(\add_83_2_C130_G3/carry[8] ), 
        .CO(\add_83_2_C130_G3/carry[9] ), .S(\tmp_A_neg[2][8] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_9  ( .A(N10), .B(\add_83_2_C130_G3/carry[9] ), 
        .CO(\add_83_2_C130_G3/carry[10] ), .S(\tmp_A_neg[2][9] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_10  ( .A(N9), .B(\add_83_2_C130_G3/carry[10] ), 
        .CO(\add_83_2_C130_G3/carry[11] ), .S(\tmp_A_neg[2][10] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_11  ( .A(N8), .B(\add_83_2_C130_G3/carry[11] ), 
        .CO(\add_83_2_C130_G3/carry[12] ), .S(\tmp_A_neg[2][11] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_12  ( .A(N7), .B(\add_83_2_C130_G3/carry[12] ), 
        .CO(\add_83_2_C130_G3/carry[13] ), .S(\tmp_A_neg[2][12] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_13  ( .A(N6), .B(\add_83_2_C130_G3/carry[13] ), 
        .CO(\add_83_2_C130_G3/carry[14] ), .S(\tmp_A_neg[2][13] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_14  ( .A(N5), .B(\add_83_2_C130_G3/carry[14] ), 
        .CO(\add_83_2_C130_G3/carry[15] ), .S(\tmp_A_neg[2][14] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_15  ( .A(N4), .B(\add_83_2_C130_G3/carry[15] ), 
        .CO(\add_83_2_C130_G3/carry[16] ), .S(\tmp_A_neg[2][15] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_16  ( .A(N3), .B(\add_83_2_C130_G3/carry[16] ), 
        .CO(\add_83_2_C130_G3/carry[17] ), .S(\tmp_A_neg[2][16] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_17  ( .A(N2), .B(\add_83_2_C130_G3/carry[17] ), 
        .CO(\add_83_2_C130_G3/carry[18] ), .S(\tmp_A_neg[2][17] ) );
  HA_X1 \add_83_2_C130_G3/U1_1_18  ( .A(N1), .B(\add_83_2_C130_G3/carry[18] ), 
        .CO(\add_83_2_C130_G3/carry[19] ), .S(\tmp_A_neg[2][18] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_4  ( .A(n53), .B(n40), .CO(
        \add_83_2_C132_G2/carry[5] ), .S(\tmp_A_neg_double[1][4] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_5  ( .A(N13), .B(\add_83_2_C132_G2/carry[5] ), 
        .CO(\add_83_2_C132_G2/carry[6] ), .S(\tmp_A_neg_double[1][5] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_6  ( .A(N12), .B(\add_83_2_C132_G2/carry[6] ), 
        .CO(\add_83_2_C132_G2/carry[7] ), .S(\tmp_A_neg_double[1][6] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_7  ( .A(N11), .B(\add_83_2_C132_G2/carry[7] ), 
        .CO(\add_83_2_C132_G2/carry[8] ), .S(\tmp_A_neg_double[1][7] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_8  ( .A(N10), .B(\add_83_2_C132_G2/carry[8] ), 
        .CO(\add_83_2_C132_G2/carry[9] ), .S(\tmp_A_neg_double[1][8] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_9  ( .A(N9), .B(\add_83_2_C132_G2/carry[9] ), 
        .CO(\add_83_2_C132_G2/carry[10] ), .S(\tmp_A_neg_double[1][9] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_10  ( .A(N8), .B(\add_83_2_C132_G2/carry[10] ), 
        .CO(\add_83_2_C132_G2/carry[11] ), .S(\tmp_A_neg_double[1][10] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_11  ( .A(N7), .B(\add_83_2_C132_G2/carry[11] ), 
        .CO(\add_83_2_C132_G2/carry[12] ), .S(\tmp_A_neg_double[1][11] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_12  ( .A(N6), .B(\add_83_2_C132_G2/carry[12] ), 
        .CO(\add_83_2_C132_G2/carry[13] ), .S(\tmp_A_neg_double[1][12] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_15  ( .A(N3), .B(n20), .CO(
        \add_83_2_C132_G2/carry[16] ), .S(\tmp_A_neg_double[1][15] ) );
  HA_X1 \add_83_2_C132_G2/U1_1_16  ( .A(N2), .B(\add_83_2_C132_G2/carry[16] ), 
        .CO(\add_83_2_C132_G2/carry[17] ), .S(\tmp_A_neg_double[1][16] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_3  ( .A(n53), .B(\add_83_2_C130_G8/carry[15] ), 
        .CO(\add_83_2_C130_G2/carry[4] ), .S(\tmp_A_neg[1][3] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_4  ( .A(N13), .B(\add_83_2_C130_G2/carry[4] ), 
        .CO(\add_83_2_C130_G2/carry[5] ), .S(\tmp_A_neg[1][4] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_5  ( .A(N12), .B(\add_83_2_C130_G2/carry[5] ), 
        .CO(\add_83_2_C130_G2/carry[6] ), .S(\tmp_A_neg[1][5] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_6  ( .A(N11), .B(\add_83_2_C130_G2/carry[6] ), 
        .CO(\add_83_2_C130_G2/carry[7] ), .S(\tmp_A_neg[1][6] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_7  ( .A(N10), .B(\add_83_2_C130_G2/carry[7] ), 
        .CO(\add_83_2_C130_G2/carry[8] ), .S(\tmp_A_neg[1][7] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_9  ( .A(N8), .B(\add_83_2_C130_G2/carry[9] ), 
        .CO(\add_83_2_C130_G2/carry[10] ), .S(\tmp_A_neg[1][9] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_10  ( .A(N7), .B(\add_83_2_C130_G2/carry[10] ), 
        .CO(\add_83_2_C130_G2/carry[11] ), .S(\tmp_A_neg[1][10] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_11  ( .A(N6), .B(\add_83_2_C130_G2/carry[11] ), 
        .CO(\add_83_2_C130_G2/carry[12] ), .S(\tmp_A_neg[1][11] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_12  ( .A(N5), .B(\add_83_2_C130_G2/carry[12] ), 
        .CO(\add_83_2_C130_G2/carry[13] ), .S(\tmp_A_neg[1][12] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_13  ( .A(N4), .B(\add_83_2_C130_G2/carry[13] ), 
        .CO(\add_83_2_C130_G2/carry[14] ), .S(\tmp_A_neg[1][13] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_14  ( .A(N3), .B(\add_83_2_C130_G2/carry[14] ), 
        .CO(\add_83_2_C130_G2/carry[15] ), .S(\tmp_A_neg[1][14] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_15  ( .A(N2), .B(\add_83_2_C130_G2/carry[15] ), 
        .CO(\add_83_2_C130_G2/carry[16] ), .S(\tmp_A_neg[1][15] ) );
  HA_X1 \add_83_2_C130_G2/U1_1_16  ( .A(N1), .B(\add_83_2_C130_G2/carry[16] ), 
        .CO(\add_83_2_C130_G2/carry[17] ), .S(\tmp_A_neg[1][16] ) );
  HA_X1 \add_83_2_C111/U1_1_5  ( .A(N11), .B(n50), .CO(
        \add_83_2_C111/carry[6] ), .S(\tmp_A_neg_double[0][5] ) );
  HA_X1 \add_83_2_C111/U1_1_6  ( .A(N10), .B(\add_83_2_C111/carry[6] ), .CO(
        \add_83_2_C111/carry[7] ), .S(\tmp_A_neg_double[0][6] ) );
  HA_X1 \add_83_2_C111/U1_1_9  ( .A(N7), .B(n49), .CO(
        \add_83_2_C111/carry[10] ), .S(\tmp_A_neg_double[0][9] ) );
  HA_X1 \add_109/U1_1_4  ( .A(N11), .B(\add_109/carry[4] ), .CO(
        \add_109/carry[5] ), .S(\tmp_A_neg[0][4] ) );
  HA_X1 \add_109/U1_1_5  ( .A(N10), .B(\add_109/carry[5] ), .CO(
        \add_109/carry[6] ), .S(\tmp_A_neg[0][5] ) );
  HA_X1 \add_109/U1_1_11  ( .A(N4), .B(n36), .CO(\add_109/carry[12] ), .S(
        \tmp_A_neg[0][11] ) );
  HA_X1 \add_109/U1_1_14  ( .A(n46), .B(N1), .CO(\add_109/carry[15] ), .S(
        \tmp_A_neg[0][14] ) );
  AND2_X4 U20 ( .A1(N7), .A2(\add_109/carry[8] ), .ZN(n18) );
  AND2_X4 U21 ( .A1(N6), .A2(n18), .ZN(n19) );
  AND2_X4 U22 ( .A1(N4), .A2(n24), .ZN(n20) );
  INV_X2 U23 ( .A(n39), .ZN(\add_109/carry[2] ) );
  NAND2_X2 U24 ( .A1(n53), .A2(n54), .ZN(n39) );
  AND2_X4 U25 ( .A1(n31), .A2(n85), .ZN(\tmp_A_neg_double[1][31] ) );
  NAND2_X2 U26 ( .A1(N1), .A2(\add_83_2_C132_G2/carry[17] ), .ZN(n31) );
  AND2_X4 U27 ( .A1(N5), .A2(\add_83_2_C132_G2/carry[13] ), .ZN(n24) );
  AND2_X4 U28 ( .A1(N9), .A2(\add_109/carry[6] ), .ZN(n25) );
  NAND2_X4 U29 ( .A1(N8), .A2(n25), .ZN(n33) );
  AND2_X2 U30 ( .A1(N9), .A2(n34), .ZN(n21) );
  INV_X2 U31 ( .A(A[6]), .ZN(N9) );
  INV_X4 U32 ( .A(n33), .ZN(\add_109/carry[8] ) );
  INV_X1 U33 ( .A(A[14]), .ZN(N1) );
  INV_X16 U34 ( .A(A[0]), .ZN(n40) );
  AND2_X1 U35 ( .A1(N12), .A2(n48), .ZN(n50) );
  AND2_X1 U36 ( .A1(N8), .A2(n21), .ZN(n49) );
  INV_X1 U37 ( .A(n43), .ZN(\add_83_2_C111/carry[16] ) );
  NAND2_X1 U38 ( .A1(N1), .A2(n23), .ZN(n43) );
  INV_X8 U39 ( .A(A[2]), .ZN(N13) );
  INV_X1 U40 ( .A(A[10]), .ZN(N5) );
  INV_X1 U41 ( .A(A[11]), .ZN(N4) );
  INV_X4 U42 ( .A(A[4]), .ZN(N11) );
  INV_X2 U43 ( .A(A[5]), .ZN(N10) );
  INV_X1 U44 ( .A(A[8]), .ZN(N7) );
  INV_X1 U45 ( .A(A[9]), .ZN(N6) );
  INV_X1 U46 ( .A(A[13]), .ZN(N2) );
  INV_X4 U47 ( .A(A[3]), .ZN(N12) );
  INV_X16 U48 ( .A(A[0]), .ZN(\add_83_2_C130_G8/carry[15] ) );
  INV_X1 U49 ( .A(A[7]), .ZN(N8) );
  BUF_X1 U50 ( .A(\tmp_A_neg[0][31] ), .Z(n52) );
  AND2_X2 U51 ( .A1(N13), .A2(\add_109/carry[2] ), .ZN(n22) );
  AND2_X1 U52 ( .A1(N2), .A2(n47), .ZN(n23) );
  AND2_X1 U53 ( .A1(N6), .A2(\add_83_2_C111/carry[10] ), .ZN(n26) );
  AND2_X1 U54 ( .A1(N5), .A2(n26), .ZN(n27) );
  INV_X16 U55 ( .A(A[1]), .ZN(n53) );
  AND2_X2 U56 ( .A1(N13), .A2(n51), .ZN(n48) );
  INV_X1 U57 ( .A(n31), .ZN(\add_83_2_C132_G2/carry[18] ) );
  INV_X2 U58 ( .A(\tmp_A_neg_double[1][31] ), .ZN(n44) );
  INV_X4 U59 ( .A(n44), .ZN(n45) );
  AND2_X4 U60 ( .A1(N3), .A2(n35), .ZN(n46) );
  AND2_X2 U61 ( .A1(\add_109/carry[12] ), .A2(N2), .ZN(n35) );
  XOR2_X1 U62 ( .A(N5), .B(\add_83_2_C132_G2/carry[13] ), .Z(
        \tmp_A_neg_double[1][13] ) );
  XOR2_X1 U63 ( .A(N12), .B(n22), .Z(\tmp_A_neg[0][3] ) );
  INV_X2 U64 ( .A(n28), .ZN(\add_109/carry[4] ) );
  NAND2_X2 U65 ( .A1(N12), .A2(n22), .ZN(n28) );
  XOR2_X1 U66 ( .A(N4), .B(n24), .Z(\tmp_A_neg_double[1][14] ) );
  AND2_X2 U67 ( .A1(n48), .A2(n30), .ZN(n29) );
  AND2_X1 U68 ( .A1(N12), .A2(N11), .ZN(n30) );
  XOR2_X1 U69 ( .A(N2), .B(n47), .Z(\tmp_A_neg_double[0][14] ) );
  XOR2_X1 U70 ( .A(N1), .B(\add_83_2_C132_G2/carry[17] ), .Z(
        \tmp_A_neg_double[1][17] ) );
  INV_X16 U71 ( .A(A[0]), .ZN(n54) );
  XOR2_X1 U72 ( .A(N9), .B(\add_109/carry[6] ), .Z(\tmp_A_neg[0][6] ) );
  XOR2_X1 U73 ( .A(N9), .B(\add_83_2_C130_G2/carry[8] ), .Z(\tmp_A_neg[1][8] )
         );
  INV_X2 U74 ( .A(n32), .ZN(\add_83_2_C130_G2/carry[9] ) );
  NAND2_X1 U75 ( .A1(N9), .A2(\add_83_2_C130_G2/carry[8] ), .ZN(n32) );
  XNOR2_X1 U76 ( .A(A[15]), .B(\add_83_2_C132_G2/carry[18] ), .ZN(
        \tmp_A_neg_double[1][18] ) );
  XOR2_X1 U77 ( .A(N6), .B(\add_83_2_C111/carry[10] ), .Z(
        \tmp_A_neg_double[0][10] ) );
  XOR2_X1 U78 ( .A(N8), .B(n25), .Z(\tmp_A_neg[0][7] ) );
  AND2_X2 U79 ( .A1(N10), .A2(n29), .ZN(n34) );
  XOR2_X1 U80 ( .A(N7), .B(\add_109/carry[8] ), .Z(\tmp_A_neg[0][8] ) );
  XOR2_X1 U81 ( .A(N9), .B(\add_83_2_C111/carry[7] ), .Z(
        \tmp_A_neg_double[0][7] ) );
  AND2_X1 U82 ( .A1(n43), .A2(n85), .ZN(\tmp_A_neg_double[0][31] ) );
  XOR2_X1 U83 ( .A(N6), .B(n18), .Z(\tmp_A_neg[0][9] ) );
  AND2_X4 U84 ( .A1(N5), .A2(n19), .ZN(n36) );
  XNOR2_X1 U85 ( .A(A[12]), .B(\add_109/carry[12] ), .ZN(\tmp_A_neg[0][12] )
         );
  XOR2_X1 U86 ( .A(N5), .B(n26), .Z(\tmp_A_neg_double[0][11] ) );
  XOR2_X1 U87 ( .A(N5), .B(n19), .Z(\tmp_A_neg[0][10] ) );
  AND2_X1 U88 ( .A1(n27), .A2(n37), .ZN(n47) );
  INV_X1 U89 ( .A(A[1]), .ZN(n41) );
  AND2_X1 U90 ( .A1(N4), .A2(N3), .ZN(n37) );
  AND2_X1 U91 ( .A1(N4), .A2(n27), .ZN(n38) );
  XOR2_X1 U92 ( .A(n41), .B(n57), .Z(\tmp_A_neg[0][1] ) );
  XOR2_X1 U93 ( .A(N4), .B(n27), .Z(\tmp_A_neg_double[0][12] ) );
  AND2_X1 U94 ( .A1(N3), .A2(\add_109/carry[12] ), .ZN(n42) );
  XOR2_X1 U95 ( .A(N1), .B(n23), .Z(\tmp_A_neg_double[0][15] ) );
  XOR2_X1 U96 ( .A(N13), .B(\add_109/carry[2] ), .Z(\tmp_A_neg[0][2] ) );
  INV_X1 U97 ( .A(A[12]), .ZN(N3) );
  NOR2_X1 U98 ( .A1(\add_83_2_C130_G3/carry[19] ), .A2(n70), .ZN(
        \tmp_A_neg[2][31] ) );
  NOR2_X1 U99 ( .A1(\add_83_2_C132_G3/carry[20] ), .A2(n70), .ZN(
        \tmp_A_neg_double[2][31] ) );
  NOR2_X1 U100 ( .A1(\add_83_2_C130_G4/carry[21] ), .A2(n70), .ZN(
        \tmp_A_neg[3][31] ) );
  INV_X1 U101 ( .A(n78), .ZN(n60) );
  INV_X1 U102 ( .A(n79), .ZN(n59) );
  INV_X1 U103 ( .A(n83), .ZN(n61) );
  INV_X1 U104 ( .A(n77), .ZN(n58) );
  INV_X1 U105 ( .A(n84), .ZN(n67) );
  NOR2_X1 U106 ( .A1(\add_83_2_C132_G4/carry[22] ), .A2(n70), .ZN(
        \tmp_A_neg_double[3][31] ) );
  INV_X1 U107 ( .A(n85), .ZN(n69) );
  INV_X1 U108 ( .A(n85), .ZN(n68) );
  AND2_X1 U109 ( .A1(n53), .A2(n40), .ZN(n51) );
  INV_X1 U110 ( .A(n83), .ZN(n62) );
  INV_X1 U111 ( .A(n84), .ZN(n63) );
  INV_X1 U112 ( .A(n83), .ZN(n64) );
  INV_X1 U113 ( .A(n84), .ZN(n65) );
  INV_X1 U114 ( .A(n85), .ZN(n66) );
  BUF_X1 U115 ( .A(A[0]), .Z(n55) );
  NOR2_X1 U116 ( .A1(\add_109/carry[15] ), .A2(n69), .ZN(\tmp_A_neg[0][31] )
         );
  INV_X1 U117 ( .A(n55), .ZN(n56) );
  NOR2_X2 U118 ( .A1(\add_83_2_C130_G2/carry[17] ), .A2(n69), .ZN(
        \tmp_A_neg[1][31] ) );
  XOR2_X1 U119 ( .A(n41), .B(n57), .Z(\tmp_A_neg_double[0][2] ) );
  XOR2_X1 U120 ( .A(N13), .B(n51), .Z(\tmp_A_neg_double[0][3] ) );
  XOR2_X1 U121 ( .A(N12), .B(n48), .Z(\tmp_A_neg_double[0][4] ) );
  XOR2_X1 U122 ( .A(N2), .B(n42), .Z(\tmp_A_neg[0][13] ) );
  XOR2_X1 U123 ( .A(N8), .B(n21), .Z(\tmp_A_neg_double[0][8] ) );
  XOR2_X1 U124 ( .A(N3), .B(n38), .Z(\tmp_A_neg_double[0][13] ) );
  INV_X1 U125 ( .A(n55), .ZN(n57) );
  INV_X1 U126 ( .A(n86), .ZN(n70) );
  INV_X1 U127 ( .A(A[15]), .ZN(n71) );
  INV_X1 U128 ( .A(A[15]), .ZN(n72) );
  INV_X1 U129 ( .A(A[15]), .ZN(n73) );
  INV_X1 U130 ( .A(A[15]), .ZN(n74) );
  INV_X1 U131 ( .A(A[15]), .ZN(n75) );
  INV_X1 U132 ( .A(A[15]), .ZN(n76) );
  INV_X1 U133 ( .A(A[15]), .ZN(n77) );
  INV_X1 U134 ( .A(A[15]), .ZN(n78) );
  INV_X1 U135 ( .A(A[15]), .ZN(n79) );
  INV_X1 U136 ( .A(A[15]), .ZN(n80) );
  INV_X1 U137 ( .A(A[15]), .ZN(n81) );
  INV_X1 U138 ( .A(A[15]), .ZN(n82) );
  INV_X1 U139 ( .A(A[15]), .ZN(n83) );
  INV_X1 U140 ( .A(A[15]), .ZN(n84) );
  INV_X1 U141 ( .A(A[15]), .ZN(n85) );
  INV_X1 U142 ( .A(A[15]), .ZN(n86) );
  XOR2_X1 U143 ( .A(n80), .B(\add_109/carry[15] ), .Z(\tmp_A_neg[0][15] ) );
  XOR2_X1 U144 ( .A(n81), .B(\add_83_2_C111/carry[16] ), .Z(
        \tmp_A_neg_double[0][16] ) );
  XOR2_X1 U145 ( .A(n80), .B(\add_83_2_C130_G2/carry[17] ), .Z(
        \tmp_A_neg[1][17] ) );
  XOR2_X1 U146 ( .A(n80), .B(\add_83_2_C130_G3/carry[19] ), .Z(
        \tmp_A_neg[2][19] ) );
  XOR2_X1 U147 ( .A(n82), .B(\add_83_2_C132_G3/carry[20] ), .Z(
        \tmp_A_neg_double[2][20] ) );
  XOR2_X1 U148 ( .A(n81), .B(\add_83_2_C130_G4/carry[21] ), .Z(
        \tmp_A_neg[3][21] ) );
  XOR2_X1 U149 ( .A(n82), .B(\add_83_2_C132_G4/carry[22] ), .Z(
        \tmp_A_neg_double[3][22] ) );
  XOR2_X1 U150 ( .A(n81), .B(\add_83_2_C130_G5/carry[23] ), .Z(
        \tmp_A_neg[4][23] ) );
  NOR2_X1 U151 ( .A1(\add_83_2_C130_G5/carry[23] ), .A2(n70), .ZN(
        \tmp_A_neg[4][31] ) );
  XOR2_X1 U152 ( .A(n82), .B(\add_83_2_C132_G5/carry[24] ), .Z(
        \tmp_A_neg_double[4][24] ) );
  NOR2_X1 U153 ( .A1(\add_83_2_C132_G5/carry[24] ), .A2(n70), .ZN(
        \tmp_A_neg_double[4][31] ) );
  XOR2_X1 U154 ( .A(\add_83_2_C130_G7/carry[31] ), .B(n77), .Z(
        \tmp_A_neg[6][31] ) );
  XOR2_X1 U155 ( .A(\add_83_2_C132_G7/carry[31] ), .B(n78), .Z(
        \tmp_A_neg_double[6][31] ) );
  XOR2_X1 U156 ( .A(\add_83_2_C130_G8/carry[31] ), .B(n78), .Z(
        \tmp_A_neg[7][31] ) );
  XOR2_X1 U157 ( .A(\add_83_2_C132_G8/carry[31] ), .B(n79), .Z(
        \tmp_A_neg_double[7][31] ) );
endmodule

