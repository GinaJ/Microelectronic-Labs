
module ND2_95 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module MUX21_GENERIC_N4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_7 UIV ( .A(SEL), .Y(SB) );
  ND2_84 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_83 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_82 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_81 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_80 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_79 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_78 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_77 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_76 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_75 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_74 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_73 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_6 UIV ( .A(SEL), .Y(SB) );
  ND2_72 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_71 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_70 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_69 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_68 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_67 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_66 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_65 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_64 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_63 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_62 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_61 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_5 UIV ( .A(SEL), .Y(SB) );
  ND2_60 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_59 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_58 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_57 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_56 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_55 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_54 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_53 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_52 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_51 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_50 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_49 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_4 UIV ( .A(SEL), .Y(SB) );
  ND2_48 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_47 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_46 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_45 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_44 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_43 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_42 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_41 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_40 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_39 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_38 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_37 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB, n1;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_3 UIV ( .A(SEL), .Y(SB) );
  ND2_36 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_35 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_34 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_33 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_32 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_31 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_30 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_29 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_28 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_27 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_26 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_25 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X2 U1 ( .A(SEL), .Z(n1) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB, n1;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_2 UIV ( .A(SEL), .Y(SB) );
  ND2_24 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_23 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_22 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_21 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_20 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_19 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_18 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_17 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_16 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_15 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_14 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_13 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X2 U1 ( .A(SEL), .Z(n1) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB, n1;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_1 UIV ( .A(SEL), .Y(SB) );
  ND2_12 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  ND2_11 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_10 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_9 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  ND2_8 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_7 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_6 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  ND2_5 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_4 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_3 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  ND2_2 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_1 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  BUF_X2 U1 ( .A(SEL), .Z(n1) );
endmodule


module RCA_generic_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module cs_generic_N4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_14 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_13 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_7 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_12 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_11 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_6 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_10 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_9 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_5 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_8 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_7 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_4 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_6 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_5 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_3 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_4 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_3 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_2 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module cs_generic_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_2 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_1 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_1 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module block_pg_26 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_25 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_24 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_23 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_22 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module block_pg_21 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_20 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_19 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_18 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_17 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_16 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_15 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_14 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_13 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_12 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module block_pg_11 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module block_pg_10 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_9 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module block_pg_8 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_7 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_6 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AND2_X1 U3 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
endmodule


module block_pg_5 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module block_pg_4 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_3 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_2 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_pg_1 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n3;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Gij) );
endmodule


module block_g_9 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Gij) );
endmodule


module block_g_8 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_g_7 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n3) );
endmodule


module block_g_6 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U2 ( .A1(Gk1j), .A2(Pik), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module block_g_5 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n3) );
endmodule


module block_g_4 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n3) );
endmodule


module block_g_3 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U2 ( .A1(Gk1j), .A2(Pik), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module block_g_2 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U2 ( .A1(Gk1j), .A2(Pik), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module block_g_1 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gik), .ZN(n2) );
  NAND2_X1 U2 ( .A1(Gk1j), .A2(Pik), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(Gij) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_GENERIC_N4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  IV_0 UIV ( .A(SEL), .Y(SB) );
  ND2_0 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  ND2_95 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  ND2_94 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  ND2_93 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  ND2_92 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  ND2_91 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  ND2_90 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  ND2_89 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  ND2_88 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  ND2_87 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  ND2_86 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  ND2_85 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
endmodule


module RCA_generic_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module cs_generic_N4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_generic_N4_0 UADDER1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_generic_N4_15 UADDER2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_0 U1 ( .A(S2), .B(S1), .SEL(Ci), .Y(S) );
endmodule


module block_pg_0 ( Pik, Pk1j, Gik, Gk1j, Pij, Gij );
  input Pik, Pk1j, Gik, Gk1j;
  output Pij, Gij;
  wire   n2;

  AND2_X1 U1 ( .A1(Pk1j), .A2(Pik), .ZN(Pij) );
  INV_X1 U2 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U3 ( .B1(Gk1j), .B2(Pik), .A(Gik), .ZN(n2) );
endmodule


module block_g_0 ( Pik, Gik, Gk1j, Gij );
  input Pik, Gik, Gk1j;
  output Gij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gij) );
  AOI21_X1 U2 ( .B1(Pik), .B2(Gk1j), .A(Gik), .ZN(n2) );
endmodule


module Sum_generator_Nbit32_Nblock8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  cs_generic_N4_0 cs_gen_1 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  cs_generic_N4_7 cs_gen_2 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  cs_generic_N4_6 cs_gen_3 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  cs_generic_N4_5 cs_gen_4 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  cs_generic_N4_4 cs_gen_5 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  cs_generic_N4_3 cs_gen_6 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  cs_generic_N4_2 cs_gen_7 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  cs_generic_N4_1 cs_gen_8 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module sparce_tree_POWER5 ( A, B, Ci, Cout );
  input [32:1] A;
  input [32:1] B;
  output [8:0] Cout;
  input Ci;
  wire   Ci, n10, n11, n12, p1, g1, \matrixG[16][16] , \matrixG[16][15] ,
         \matrixG[16][13] , \matrixG[16][9] , \matrixG[15][15] ,
         \matrixG[14][14] , \matrixG[14][13] , \matrixG[13][13] ,
         \matrixG[12][12] , \matrixG[12][11] , \matrixG[12][9] ,
         \matrixG[11][11] , \matrixG[10][10] , \matrixG[10][9] ,
         \matrixG[9][9] , \matrixG[8][8] , \matrixG[8][7] , \matrixG[8][5] ,
         \matrixG[7][7] , \matrixG[6][6] , \matrixG[6][5] , \matrixG[5][5] ,
         \matrixG[4][4] , \matrixG[4][3] , \matrixG[3][3] , \matrixG[2][2] ,
         \matrixG[2][1] , \matrixG[1][1] , \matrixP[16][16] ,
         \matrixP[16][15] , \matrixP[16][13] , \matrixP[16][9] ,
         \matrixP[15][15] , \matrixP[14][14] , \matrixP[14][13] ,
         \matrixP[13][13] , \matrixP[12][12] , \matrixP[12][11] ,
         \matrixP[12][9] , \matrixP[11][11] , \matrixP[10][10] ,
         \matrixP[10][9] , \matrixP[9][9] , \matrixP[8][8] , \matrixP[8][7] ,
         \matrixP[8][5] , \matrixP[7][7] , \matrixP[6][6] , \matrixP[6][5] ,
         \matrixP[5][5] , \matrixP[4][4] , \matrixP[4][3] , \matrixP[3][3] ,
         \matrixP[2][2] , \matrixP[32][32] , \matrixP[32][31] ,
         \matrixP[32][29] , \matrixP[32][25] , \matrixP[32][17] ,
         \matrixP[31][31] , \matrixP[30][30] , \matrixP[30][29] ,
         \matrixP[29][29] , \matrixP[28][28] , \matrixP[28][27] ,
         \matrixP[28][25] , \matrixP[28][17] , \matrixP[27][27] ,
         \matrixP[26][26] , \matrixP[26][25] , \matrixP[25][25] ,
         \matrixP[24][24] , \matrixP[24][23] , \matrixP[24][21] ,
         \matrixP[24][17] , \matrixP[23][23] , \matrixP[22][22] ,
         \matrixP[22][21] , \matrixP[21][21] , \matrixP[20][20] ,
         \matrixP[20][19] , \matrixP[20][17] , \matrixP[19][19] ,
         \matrixP[18][18] , \matrixP[18][17] , \matrixP[17][17] ,
         \matrixG[32][32] , \matrixG[32][31] , \matrixG[32][29] ,
         \matrixG[32][25] , \matrixG[32][17] , \matrixG[31][31] ,
         \matrixG[30][30] , \matrixG[30][29] , \matrixG[29][29] ,
         \matrixG[28][28] , \matrixG[28][27] , \matrixG[28][25] ,
         \matrixG[28][17] , \matrixG[27][27] , \matrixG[26][26] ,
         \matrixG[26][25] , \matrixG[25][25] , \matrixG[24][24] ,
         \matrixG[24][23] , \matrixG[24][21] , \matrixG[24][17] ,
         \matrixG[23][23] , \matrixG[22][22] , \matrixG[22][21] ,
         \matrixG[21][21] , \matrixG[20][20] , \matrixG[20][19] ,
         \matrixG[20][17] , \matrixG[19][19] , \matrixG[18][18] ,
         \matrixG[18][17] , \matrixG[17][17] , n1, n2, n3, n4, n5, n8;
  assign Cout[0] = Ci;

  block_g_0 blkg_Cin_0 ( .Pik(p1), .Gik(g1), .Gk1j(Ci), .Gij(\matrixG[1][1] )
         );
  block_g_9 blkg_1_1 ( .Pik(\matrixP[2][2] ), .Gik(\matrixG[2][2] ), .Gk1j(
        \matrixG[1][1] ), .Gij(\matrixG[2][1] ) );
  block_pg_0 blkpg_1_2 ( .Pik(\matrixP[4][4] ), .Pk1j(\matrixP[3][3] ), .Gik(
        \matrixG[4][4] ), .Gk1j(\matrixG[3][3] ), .Pij(\matrixP[4][3] ), .Gij(
        \matrixG[4][3] ) );
  block_pg_26 blkpg_1_3 ( .Pik(\matrixP[6][6] ), .Pk1j(\matrixP[5][5] ), .Gik(
        \matrixG[6][6] ), .Gk1j(\matrixG[5][5] ), .Pij(\matrixP[6][5] ), .Gij(
        \matrixG[6][5] ) );
  block_pg_25 blkpg_1_4 ( .Pik(\matrixP[8][8] ), .Pk1j(\matrixP[7][7] ), .Gik(
        \matrixG[8][8] ), .Gk1j(\matrixG[7][7] ), .Pij(\matrixP[8][7] ), .Gij(
        \matrixG[8][7] ) );
  block_pg_24 blkpg_1_5 ( .Pik(\matrixP[10][10] ), .Pk1j(\matrixP[9][9] ), 
        .Gik(\matrixG[10][10] ), .Gk1j(\matrixG[9][9] ), .Pij(\matrixP[10][9] ), .Gij(\matrixG[10][9] ) );
  block_pg_23 blkpg_1_6 ( .Pik(\matrixP[12][12] ), .Pk1j(\matrixP[11][11] ), 
        .Gik(\matrixG[12][12] ), .Gk1j(\matrixG[11][11] ), .Pij(
        \matrixP[12][11] ), .Gij(\matrixG[12][11] ) );
  block_pg_22 blkpg_1_7 ( .Pik(\matrixP[14][14] ), .Pk1j(\matrixP[13][13] ), 
        .Gik(\matrixG[14][14] ), .Gk1j(\matrixG[13][13] ), .Pij(
        \matrixP[14][13] ), .Gij(\matrixG[14][13] ) );
  block_pg_21 blkpg_1_8 ( .Pik(\matrixP[16][16] ), .Pk1j(\matrixP[15][15] ), 
        .Gik(\matrixG[16][16] ), .Gk1j(\matrixG[15][15] ), .Pij(
        \matrixP[16][15] ), .Gij(\matrixG[16][15] ) );
  block_pg_20 blkpg_1_9 ( .Pik(\matrixP[18][18] ), .Pk1j(\matrixP[17][17] ), 
        .Gik(\matrixG[18][18] ), .Gk1j(\matrixG[17][17] ), .Pij(
        \matrixP[18][17] ), .Gij(\matrixG[18][17] ) );
  block_pg_19 blkpg_1_10 ( .Pik(\matrixP[20][20] ), .Pk1j(\matrixP[19][19] ), 
        .Gik(\matrixG[20][20] ), .Gk1j(\matrixG[19][19] ), .Pij(
        \matrixP[20][19] ), .Gij(\matrixG[20][19] ) );
  block_pg_18 blkpg_1_11 ( .Pik(\matrixP[22][22] ), .Pk1j(\matrixP[21][21] ), 
        .Gik(\matrixG[22][22] ), .Gk1j(\matrixG[21][21] ), .Pij(
        \matrixP[22][21] ), .Gij(\matrixG[22][21] ) );
  block_pg_17 blkpg_1_12 ( .Pik(\matrixP[24][24] ), .Pk1j(\matrixP[23][23] ), 
        .Gik(\matrixG[24][24] ), .Gk1j(\matrixG[23][23] ), .Pij(
        \matrixP[24][23] ), .Gij(\matrixG[24][23] ) );
  block_pg_16 blkpg_1_13 ( .Pik(\matrixP[26][26] ), .Pk1j(\matrixP[25][25] ), 
        .Gik(\matrixG[26][26] ), .Gk1j(\matrixG[25][25] ), .Pij(
        \matrixP[26][25] ), .Gij(\matrixG[26][25] ) );
  block_pg_15 blkpg_1_14 ( .Pik(\matrixP[28][28] ), .Pk1j(\matrixP[27][27] ), 
        .Gik(\matrixG[28][28] ), .Gk1j(\matrixG[27][27] ), .Pij(
        \matrixP[28][27] ), .Gij(\matrixG[28][27] ) );
  block_pg_14 blkpg_1_15 ( .Pik(\matrixP[30][30] ), .Pk1j(\matrixP[29][29] ), 
        .Gik(\matrixG[30][30] ), .Gk1j(\matrixG[29][29] ), .Pij(
        \matrixP[30][29] ), .Gij(\matrixG[30][29] ) );
  block_pg_13 blkpg_1_16 ( .Pik(\matrixP[32][32] ), .Pk1j(\matrixP[31][31] ), 
        .Gik(\matrixG[32][32] ), .Gk1j(\matrixG[31][31] ), .Pij(
        \matrixP[32][31] ), .Gij(\matrixG[32][31] ) );
  block_g_8 blkg_2_1 ( .Pik(\matrixP[4][3] ), .Gik(\matrixG[4][3] ), .Gk1j(
        \matrixG[2][1] ), .Gij(n12) );
  block_pg_12 blkpg_2_2 ( .Pik(\matrixP[8][7] ), .Pk1j(\matrixP[6][5] ), .Gik(
        \matrixG[8][7] ), .Gk1j(\matrixG[6][5] ), .Pij(\matrixP[8][5] ), .Gij(
        \matrixG[8][5] ) );
  block_pg_11 blkpg_2_3 ( .Pik(\matrixP[12][11] ), .Pk1j(\matrixP[10][9] ), 
        .Gik(\matrixG[12][11] ), .Gk1j(\matrixG[10][9] ), .Pij(
        \matrixP[12][9] ), .Gij(\matrixG[12][9] ) );
  block_pg_10 blkpg_2_4 ( .Pik(\matrixP[16][15] ), .Pk1j(\matrixP[14][13] ), 
        .Gik(\matrixG[16][15] ), .Gk1j(\matrixG[14][13] ), .Pij(
        \matrixP[16][13] ), .Gij(\matrixG[16][13] ) );
  block_pg_9 blkpg_2_5 ( .Pik(\matrixP[20][19] ), .Pk1j(\matrixP[18][17] ), 
        .Gik(\matrixG[20][19] ), .Gk1j(\matrixG[18][17] ), .Pij(
        \matrixP[20][17] ), .Gij(\matrixG[20][17] ) );
  block_pg_8 blkpg_2_6 ( .Pik(\matrixP[24][23] ), .Pk1j(\matrixP[22][21] ), 
        .Gik(\matrixG[24][23] ), .Gk1j(\matrixG[22][21] ), .Pij(
        \matrixP[24][21] ), .Gij(\matrixG[24][21] ) );
  block_pg_7 blkpg_2_7 ( .Pik(\matrixP[28][27] ), .Pk1j(\matrixP[26][25] ), 
        .Gik(\matrixG[28][27] ), .Gk1j(\matrixG[26][25] ), .Pij(
        \matrixP[28][25] ), .Gij(\matrixG[28][25] ) );
  block_pg_6 blkpg_2_8 ( .Pik(\matrixP[32][31] ), .Pk1j(\matrixP[30][29] ), 
        .Gik(\matrixG[32][31] ), .Gk1j(\matrixG[30][29] ), .Pij(
        \matrixP[32][29] ), .Gij(\matrixG[32][29] ) );
  block_g_7 blkg_3_1 ( .Pik(\matrixP[8][5] ), .Gik(\matrixG[8][5] ), .Gk1j(n12), .Gij(n11) );
  block_pg_5 blkpg_3_2 ( .Pik(\matrixP[16][13] ), .Pk1j(\matrixP[12][9] ), 
        .Gik(\matrixG[16][13] ), .Gk1j(\matrixG[12][9] ), .Pij(
        \matrixP[16][9] ), .Gij(\matrixG[16][9] ) );
  block_pg_4 blkpg_3_3 ( .Pik(\matrixP[24][21] ), .Pk1j(\matrixP[20][17] ), 
        .Gik(\matrixG[24][21] ), .Gk1j(\matrixG[20][17] ), .Pij(
        \matrixP[24][17] ), .Gij(\matrixG[24][17] ) );
  block_pg_3 blkpg_3_4 ( .Pik(\matrixP[32][29] ), .Pk1j(\matrixP[28][25] ), 
        .Gik(\matrixG[32][29] ), .Gk1j(\matrixG[28][25] ), .Pij(
        \matrixP[32][25] ), .Gij(\matrixG[32][25] ) );
  block_g_6 blkg_4_1_0 ( .Pik(\matrixP[16][9] ), .Gik(\matrixG[16][9] ), 
        .Gk1j(n11), .Gij(n10) );
  block_g_5 blkg_4_1_1 ( .Pik(\matrixP[12][9] ), .Gik(\matrixG[12][9] ), 
        .Gk1j(n1), .Gij(Cout[3]) );
  block_pg_2 blkpg_4_2_0 ( .Pik(\matrixP[32][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[32][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[32][17] ), .Gij(\matrixG[32][17] ) );
  block_pg_1 blkpg_4_2_1 ( .Pik(\matrixP[28][25] ), .Pk1j(\matrixP[24][17] ), 
        .Gik(\matrixG[28][25] ), .Gk1j(\matrixG[24][17] ), .Pij(
        \matrixP[28][17] ), .Gij(\matrixG[28][17] ) );
  block_g_4 blkg_5_1_0 ( .Pik(\matrixP[32][17] ), .Gik(\matrixG[32][17] ), 
        .Gk1j(Cout[4]), .Gij(Cout[8]) );
  block_g_3 blkg_5_1_1 ( .Pik(\matrixP[28][17] ), .Gik(\matrixG[28][17] ), 
        .Gk1j(n10), .Gij(Cout[7]) );
  block_g_2 blkg_5_1_2 ( .Pik(\matrixP[24][17] ), .Gik(\matrixG[24][17] ), 
        .Gk1j(n10), .Gij(Cout[6]) );
  block_g_1 blkg_5_1_3 ( .Pik(\matrixP[20][17] ), .Gik(\matrixG[20][17] ), 
        .Gk1j(n10), .Gij(Cout[5]) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(\matrixP[9][9] ) );
  XOR2_X1 U35 ( .A(B[8]), .B(A[8]), .Z(\matrixP[8][8] ) );
  XOR2_X1 U36 ( .A(B[7]), .B(A[7]), .Z(\matrixP[7][7] ) );
  XOR2_X1 U37 ( .A(B[6]), .B(A[6]), .Z(\matrixP[6][6] ) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(\matrixP[5][5] ) );
  XOR2_X1 U39 ( .A(B[4]), .B(A[4]), .Z(\matrixP[4][4] ) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(\matrixP[3][3] ) );
  XOR2_X1 U41 ( .A(B[32]), .B(A[32]), .Z(\matrixP[32][32] ) );
  XOR2_X1 U42 ( .A(B[31]), .B(A[31]), .Z(\matrixP[31][31] ) );
  XOR2_X1 U43 ( .A(B[30]), .B(A[30]), .Z(\matrixP[30][30] ) );
  XOR2_X1 U44 ( .A(B[2]), .B(A[2]), .Z(\matrixP[2][2] ) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(\matrixP[29][29] ) );
  XOR2_X1 U46 ( .A(B[28]), .B(A[28]), .Z(\matrixP[28][28] ) );
  XOR2_X1 U47 ( .A(B[27]), .B(A[27]), .Z(\matrixP[27][27] ) );
  XOR2_X1 U48 ( .A(B[26]), .B(A[26]), .Z(\matrixP[26][26] ) );
  XOR2_X1 U49 ( .A(B[25]), .B(A[25]), .Z(\matrixP[25][25] ) );
  XOR2_X1 U50 ( .A(B[24]), .B(A[24]), .Z(\matrixP[24][24] ) );
  XOR2_X1 U51 ( .A(B[23]), .B(A[23]), .Z(\matrixP[23][23] ) );
  XOR2_X1 U52 ( .A(B[22]), .B(A[22]), .Z(\matrixP[22][22] ) );
  XOR2_X1 U53 ( .A(B[21]), .B(A[21]), .Z(\matrixP[21][21] ) );
  XOR2_X1 U54 ( .A(B[20]), .B(A[20]), .Z(\matrixP[20][20] ) );
  XOR2_X1 U55 ( .A(B[19]), .B(A[19]), .Z(\matrixP[19][19] ) );
  XOR2_X1 U56 ( .A(B[18]), .B(A[18]), .Z(\matrixP[18][18] ) );
  XOR2_X1 U57 ( .A(B[17]), .B(A[17]), .Z(\matrixP[17][17] ) );
  XOR2_X1 U58 ( .A(B[16]), .B(A[16]), .Z(\matrixP[16][16] ) );
  XOR2_X1 U59 ( .A(B[15]), .B(A[15]), .Z(\matrixP[15][15] ) );
  XOR2_X1 U60 ( .A(B[14]), .B(A[14]), .Z(\matrixP[14][14] ) );
  XOR2_X1 U61 ( .A(B[13]), .B(A[13]), .Z(\matrixP[13][13] ) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(\matrixP[12][12] ) );
  XOR2_X1 U63 ( .A(B[11]), .B(A[11]), .Z(\matrixP[11][11] ) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(\matrixP[10][10] ) );
  BUF_X1 U1 ( .A(n11), .Z(n1) );
  BUF_X1 U2 ( .A(n10), .Z(Cout[4]) );
  AND2_X1 U3 ( .A1(B[15]), .A2(A[15]), .ZN(\matrixG[15][15] ) );
  AND2_X1 U4 ( .A1(B[16]), .A2(A[16]), .ZN(\matrixG[16][16] ) );
  AND2_X1 U5 ( .A1(B[11]), .A2(A[11]), .ZN(\matrixG[11][11] ) );
  AND2_X1 U6 ( .A1(B[12]), .A2(A[12]), .ZN(\matrixG[12][12] ) );
  AND2_X1 U7 ( .A1(B[3]), .A2(A[3]), .ZN(\matrixG[3][3] ) );
  AND2_X1 U8 ( .A1(B[4]), .A2(A[4]), .ZN(\matrixG[4][4] ) );
  AND2_X1 U9 ( .A1(B[27]), .A2(A[27]), .ZN(\matrixG[27][27] ) );
  AND2_X1 U10 ( .A1(B[28]), .A2(A[28]), .ZN(\matrixG[28][28] ) );
  AND2_X1 U11 ( .A1(B[25]), .A2(A[25]), .ZN(\matrixG[25][25] ) );
  AND2_X1 U12 ( .A1(B[26]), .A2(A[26]), .ZN(\matrixG[26][26] ) );
  AND2_X1 U13 ( .A1(B[31]), .A2(A[31]), .ZN(\matrixG[31][31] ) );
  AND2_X1 U14 ( .A1(B[32]), .A2(A[32]), .ZN(\matrixG[32][32] ) );
  AND2_X1 U15 ( .A1(B[19]), .A2(A[19]), .ZN(\matrixG[19][19] ) );
  AND2_X1 U16 ( .A1(B[20]), .A2(A[20]), .ZN(\matrixG[20][20] ) );
  AND2_X1 U17 ( .A1(B[17]), .A2(A[17]), .ZN(\matrixG[17][17] ) );
  AND2_X1 U18 ( .A1(B[18]), .A2(A[18]), .ZN(\matrixG[18][18] ) );
  AND2_X1 U19 ( .A1(B[5]), .A2(A[5]), .ZN(\matrixG[5][5] ) );
  AND2_X1 U20 ( .A1(B[6]), .A2(A[6]), .ZN(\matrixG[6][6] ) );
  AND2_X1 U21 ( .A1(B[9]), .A2(A[9]), .ZN(\matrixG[9][9] ) );
  AND2_X1 U22 ( .A1(B[10]), .A2(A[10]), .ZN(\matrixG[10][10] ) );
  AND2_X1 U23 ( .A1(B[13]), .A2(A[13]), .ZN(\matrixG[13][13] ) );
  AND2_X1 U24 ( .A1(B[14]), .A2(A[14]), .ZN(\matrixG[14][14] ) );
  AND2_X1 U25 ( .A1(B[23]), .A2(A[23]), .ZN(\matrixG[23][23] ) );
  AND2_X1 U26 ( .A1(B[24]), .A2(A[24]), .ZN(\matrixG[24][24] ) );
  AND2_X1 U27 ( .A1(B[30]), .A2(A[30]), .ZN(\matrixG[30][30] ) );
  AND2_X1 U28 ( .A1(B[29]), .A2(A[29]), .ZN(\matrixG[29][29] ) );
  AND2_X1 U29 ( .A1(B[21]), .A2(A[21]), .ZN(\matrixG[21][21] ) );
  AND2_X1 U30 ( .A1(B[22]), .A2(A[22]), .ZN(\matrixG[22][22] ) );
  AND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(\matrixG[2][2] ) );
  AND2_X1 U32 ( .A1(B[7]), .A2(A[7]), .ZN(\matrixG[7][7] ) );
  AND2_X1 U33 ( .A1(B[8]), .A2(A[8]), .ZN(\matrixG[8][8] ) );
  AND2_X1 U65 ( .A1(B[1]), .A2(A[1]), .ZN(g1) );
  NAND2_X1 U66 ( .A1(n3), .A2(B[1]), .ZN(n4) );
  NAND2_X1 U67 ( .A1(n2), .A2(A[1]), .ZN(n5) );
  NAND2_X1 U68 ( .A1(n4), .A2(n5), .ZN(p1) );
  INV_X1 U69 ( .A(B[1]), .ZN(n2) );
  INV_X1 U70 ( .A(A[1]), .ZN(n3) );
  CLKBUF_X1 U71 ( .A(n12), .Z(Cout[1]) );
  INV_X1 U72 ( .A(n1), .ZN(n8) );
  INV_X1 U73 ( .A(n8), .ZN(Cout[2]) );
endmodule


module P4adder ( A, B, Ci, S, Overf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Overf;
  wire   n1, n2;
  wire   [7:0] sCout;

  sparce_tree_POWER5 Usparce_tree ( .A(A), .B(B), .Ci(Ci), .Cout({Overf, sCout}) );
  Sum_generator_Nbit32_Nblock8 USum_generator ( .A({A[31:1], n1}), .B({B[31:1], 
        n2}), .Ci(sCout), .S(S) );
  BUF_X1 U1 ( .A(B[0]), .Z(n2) );
  BUF_X1 U2 ( .A(A[0]), .Z(n1) );
endmodule

